module FrogSpriteBram (
    input wire clk,                     // Clock signal
    input wire [4:0] sprite_x,          // X coordinate within the frog sprite (0-31)
    input wire [4:0] sprite_y,          // Y coordinate within the frog sprite (0-31)
    input wire [1:0] direction,         // Direction input: 00 = up, 01 = down, 10 = left, 11 = right
    output reg [5:0] pixel_data         // 6-bit pixel data (RGB 2-2-2)
);

    // Declare a 4096x6 bit Block RAM (BRAM) to store 32x32 frog sprites for 4 directions (up, down, left, right)
    reg [4:0] frog_bram [0:4095];       // 4096 addresses (1024 per sprite)

    // Initialize the frog sprite data for all directions
    initial begin
        /// Add more initialization here for the up-facing sprite (0 - 1023)
frog_bram[0] = 6'b000000;
frog_bram[1] = 6'b000000;
frog_bram[2] = 6'b000000;
frog_bram[3] = 6'b000000;
frog_bram[4] = 6'b000000;
frog_bram[5] = 6'b000000;
frog_bram[6] = 6'b000000;
frog_bram[7] = 6'b000000;
frog_bram[8] = 6'b000000;
frog_bram[9] = 6'b000000;
frog_bram[10] = 6'b000000;
frog_bram[11] = 6'b000000;
frog_bram[12] = 6'b000000;
frog_bram[13] = 6'b000000;
frog_bram[14] = 6'b000000;
frog_bram[15] = 6'b000000;
frog_bram[16] = 6'b000000;
frog_bram[17] = 6'b000000;
frog_bram[18] = 6'b000000;
frog_bram[19] = 6'b000000;
frog_bram[20] = 6'b000000;
frog_bram[21] = 6'b000000;
frog_bram[22] = 6'b000000;
frog_bram[23] = 6'b000000;
frog_bram[24] = 6'b000000;
frog_bram[25] = 6'b000000;
frog_bram[26] = 6'b000000;
frog_bram[27] = 6'b000000;
frog_bram[28] = 6'b000000;
frog_bram[29] = 6'b000000;
frog_bram[30] = 6'b000000;
frog_bram[31] = 6'b000000;
frog_bram[32] = 6'b000000;
frog_bram[33] = 6'b000000;
frog_bram[34] = 6'b000000;
frog_bram[35] = 6'b000000;
frog_bram[36] = 6'b000000;
frog_bram[37] = 6'b000000;
frog_bram[38] = 6'b000000;
frog_bram[39] = 6'b000000;
frog_bram[40] = 6'b000000;
frog_bram[41] = 6'b000000;
frog_bram[42] = 6'b000000;
frog_bram[43] = 6'b000000;
frog_bram[44] = 6'b000000;
frog_bram[45] = 6'b000000;
frog_bram[46] = 6'b000000;
frog_bram[47] = 6'b000000;
frog_bram[48] = 6'b000000;
frog_bram[49] = 6'b000000;
frog_bram[50] = 6'b000000;
frog_bram[51] = 6'b000000;
frog_bram[52] = 6'b000000;
frog_bram[53] = 6'b000000;
frog_bram[54] = 6'b000000;
frog_bram[55] = 6'b000000;
frog_bram[56] = 6'b000000;
frog_bram[57] = 6'b000000;
frog_bram[58] = 6'b000000;
frog_bram[59] = 6'b000000;
frog_bram[60] = 6'b000000;
frog_bram[61] = 6'b000000;
frog_bram[62] = 6'b000000;
frog_bram[63] = 6'b000000;
frog_bram[64] = 6'b000000;
frog_bram[65] = 6'b000000;
frog_bram[66] = 6'b000000;
frog_bram[67] = 6'b000000;
frog_bram[68] = 6'b000000;
frog_bram[69] = 6'b000000;
frog_bram[70] = 6'b000000;
frog_bram[71] = 6'b000000;
frog_bram[72] = 6'b000000;
frog_bram[73] = 6'b000000;
frog_bram[74] = 6'b000000;
frog_bram[75] = 6'b000000;
frog_bram[76] = 6'b000000;
frog_bram[77] = 6'b001000;
frog_bram[78] = 6'b001000;
frog_bram[79] = 6'b001100;
frog_bram[80] = 6'b001100;
frog_bram[81] = 6'b001000;
frog_bram[82] = 6'b001000;
frog_bram[83] = 6'b000000;
frog_bram[84] = 6'b000000;
frog_bram[85] = 6'b000000;
frog_bram[86] = 6'b000000;
frog_bram[87] = 6'b000000;
frog_bram[88] = 6'b000000;
frog_bram[89] = 6'b000000;
frog_bram[90] = 6'b000000;
frog_bram[91] = 6'b000000;
frog_bram[92] = 6'b000000;
frog_bram[93] = 6'b000000;
frog_bram[94] = 6'b000000;
frog_bram[95] = 6'b000000;
frog_bram[96] = 6'b000000;
frog_bram[97] = 6'b000000;
frog_bram[98] = 6'b000000;
frog_bram[99] = 6'b001100;
frog_bram[100] = 6'b001000;
frog_bram[101] = 6'b000000;
frog_bram[102] = 6'b001000;
frog_bram[103] = 6'b001000;
frog_bram[104] = 6'b000000;
frog_bram[105] = 6'b000000;
frog_bram[106] = 6'b000000;
frog_bram[107] = 6'b000000;
frog_bram[108] = 6'b001100;
frog_bram[109] = 6'b001100;
frog_bram[110] = 6'b000100;
frog_bram[111] = 6'b001100;
frog_bram[112] = 6'b001100;
frog_bram[113] = 6'b000100;
frog_bram[114] = 6'b001100;
frog_bram[115] = 6'b001100;
frog_bram[116] = 6'b000000;
frog_bram[117] = 6'b000000;
frog_bram[118] = 6'b000000;
frog_bram[119] = 6'b000000;
frog_bram[120] = 6'b001000;
frog_bram[121] = 6'b001000;
frog_bram[122] = 6'b000000;
frog_bram[123] = 6'b001000;
frog_bram[124] = 6'b001100;
frog_bram[125] = 6'b000000;
frog_bram[126] = 6'b000000;
frog_bram[127] = 6'b000000;
frog_bram[128] = 6'b000000;
frog_bram[129] = 6'b000000;
frog_bram[130] = 6'b000000;
frog_bram[131] = 6'b001100;
frog_bram[132] = 6'b001000;
frog_bram[133] = 6'b000000;
frog_bram[134] = 6'b001100;
frog_bram[135] = 6'b001000;
frog_bram[136] = 6'b000000;
frog_bram[137] = 6'b000000;
frog_bram[138] = 6'b000000;
frog_bram[139] = 6'b001000;
frog_bram[140] = 6'b001100;
frog_bram[141] = 6'b001100;
frog_bram[142] = 6'b001100;
frog_bram[143] = 6'b001100;
frog_bram[144] = 6'b001100;
frog_bram[145] = 6'b001100;
frog_bram[146] = 6'b001100;
frog_bram[147] = 6'b001100;
frog_bram[148] = 6'b001000;
frog_bram[149] = 6'b000000;
frog_bram[150] = 6'b000000;
frog_bram[151] = 6'b000000;
frog_bram[152] = 6'b001000;
frog_bram[153] = 6'b001100;
frog_bram[154] = 6'b000000;
frog_bram[155] = 6'b001000;
frog_bram[156] = 6'b001100;
frog_bram[157] = 6'b000000;
frog_bram[158] = 6'b000000;
frog_bram[159] = 6'b000000;
frog_bram[160] = 6'b000000;
frog_bram[161] = 6'b000000;
frog_bram[162] = 6'b000000;
frog_bram[163] = 6'b001100;
frog_bram[164] = 6'b000100;
frog_bram[165] = 6'b001100;
frog_bram[166] = 6'b001100;
frog_bram[167] = 6'b000000;
frog_bram[168] = 6'b000000;
frog_bram[169] = 6'b000000;
frog_bram[170] = 6'b001000;
frog_bram[171] = 6'b001000;
frog_bram[172] = 6'b001000;
frog_bram[173] = 6'b001100;
frog_bram[174] = 6'b001100;
frog_bram[175] = 6'b001100;
frog_bram[176] = 6'b001100;
frog_bram[177] = 6'b001100;
frog_bram[178] = 6'b001100;
frog_bram[179] = 6'b001100;
frog_bram[180] = 6'b001100;
frog_bram[181] = 6'b001000;
frog_bram[182] = 6'b000000;
frog_bram[183] = 6'b000000;
frog_bram[184] = 6'b000000;
frog_bram[185] = 6'b001100;
frog_bram[186] = 6'b001100;
frog_bram[187] = 6'b000100;
frog_bram[188] = 6'b001100;
frog_bram[189] = 6'b000000;
frog_bram[190] = 6'b000000;
frog_bram[191] = 6'b000000;
frog_bram[192] = 6'b000000;
frog_bram[193] = 6'b000000;
frog_bram[194] = 6'b000000;
frog_bram[195] = 6'b001100;
frog_bram[196] = 6'b001000;
frog_bram[197] = 6'b001000;
frog_bram[198] = 6'b000000;
frog_bram[199] = 6'b000000;
frog_bram[200] = 6'b000000;
frog_bram[201] = 6'b001000;
frog_bram[202] = 6'b001000;
frog_bram[203] = 6'b110000;
frog_bram[204] = 6'b110000;
frog_bram[205] = 6'b001000;
frog_bram[206] = 6'b001100;
frog_bram[207] = 6'b001100;
frog_bram[208] = 6'b001100;
frog_bram[209] = 6'b001100;
frog_bram[210] = 6'b001100;
frog_bram[211] = 6'b110000;
frog_bram[212] = 6'b110000;
frog_bram[213] = 6'b001100;
frog_bram[214] = 6'b001100;
frog_bram[215] = 6'b000000;
frog_bram[216] = 6'b000000;
frog_bram[217] = 6'b000000;
frog_bram[218] = 6'b001000;
frog_bram[219] = 6'b001000;
frog_bram[220] = 6'b001100;
frog_bram[221] = 6'b000000;
frog_bram[222] = 6'b000000;
frog_bram[223] = 6'b000000;
frog_bram[224] = 6'b000000;
frog_bram[225] = 6'b000000;
frog_bram[226] = 6'b001100;
frog_bram[227] = 6'b001100;
frog_bram[228] = 6'b001100;
frog_bram[229] = 6'b000100;
frog_bram[230] = 6'b001000;
frog_bram[231] = 6'b000000;
frog_bram[232] = 6'b000000;
frog_bram[233] = 6'b001000;
frog_bram[234] = 6'b110000;
frog_bram[235] = 6'b010000;
frog_bram[236] = 6'b010000;
frog_bram[237] = 6'b110000;
frog_bram[238] = 6'b001000;
frog_bram[239] = 6'b001100;
frog_bram[240] = 6'b001100;
frog_bram[241] = 6'b001100;
frog_bram[242] = 6'b110000;
frog_bram[243] = 6'b010000;
frog_bram[244] = 6'b010000;
frog_bram[245] = 6'b110000;
frog_bram[246] = 6'b001100;
frog_bram[247] = 6'b001100;
frog_bram[248] = 6'b000000;
frog_bram[249] = 6'b000100;
frog_bram[250] = 6'b000100;
frog_bram[251] = 6'b001100;
frog_bram[252] = 6'b001100;
frog_bram[253] = 6'b001100;
frog_bram[254] = 6'b000000;
frog_bram[255] = 6'b000000;
frog_bram[256] = 6'b000000;
frog_bram[257] = 6'b000000;
frog_bram[258] = 6'b001100;
frog_bram[259] = 6'b001100;
frog_bram[260] = 6'b001100;
frog_bram[261] = 6'b001100;
frog_bram[262] = 6'b001000;
frog_bram[263] = 6'b000000;
frog_bram[264] = 6'b001000;
frog_bram[265] = 6'b001000;
frog_bram[266] = 6'b100000;
frog_bram[267] = 6'b010000;
frog_bram[268] = 6'b010000;
frog_bram[269] = 6'b110000;
frog_bram[270] = 6'b001000;
frog_bram[271] = 6'b001100;
frog_bram[272] = 6'b001100;
frog_bram[273] = 6'b001100;
frog_bram[274] = 6'b110000;
frog_bram[275] = 6'b010000;
frog_bram[276] = 6'b010000;
frog_bram[277] = 6'b110000;
frog_bram[278] = 6'b001100;
frog_bram[279] = 6'b001100;
frog_bram[280] = 6'b000000;
frog_bram[281] = 6'b001000;
frog_bram[282] = 6'b001100;
frog_bram[283] = 6'b001100;
frog_bram[284] = 6'b001100;
frog_bram[285] = 6'b001100;
frog_bram[286] = 6'b000000;
frog_bram[287] = 6'b000000;
frog_bram[288] = 6'b000000;
frog_bram[289] = 6'b000000;
frog_bram[290] = 6'b001100;
frog_bram[291] = 6'b001100;
frog_bram[292] = 6'b001100;
frog_bram[293] = 6'b001100;
frog_bram[294] = 6'b000000;
frog_bram[295] = 6'b000000;
frog_bram[296] = 6'b001100;
frog_bram[297] = 6'b001100;
frog_bram[298] = 6'b001000;
frog_bram[299] = 6'b110000;
frog_bram[300] = 6'b110000;
frog_bram[301] = 6'b001000;
frog_bram[302] = 6'b001000;
frog_bram[303] = 6'b001100;
frog_bram[304] = 6'b001100;
frog_bram[305] = 6'b001100;
frog_bram[306] = 6'b001100;
frog_bram[307] = 6'b110000;
frog_bram[308] = 6'b110000;
frog_bram[309] = 6'b001100;
frog_bram[310] = 6'b001100;
frog_bram[311] = 6'b001100;
frog_bram[312] = 6'b000000;
frog_bram[313] = 6'b000000;
frog_bram[314] = 6'b001100;
frog_bram[315] = 6'b001100;
frog_bram[316] = 6'b001100;
frog_bram[317] = 6'b001100;
frog_bram[318] = 6'b000000;
frog_bram[319] = 6'b000000;
frog_bram[320] = 6'b000000;
frog_bram[321] = 6'b000000;
frog_bram[322] = 6'b001100;
frog_bram[323] = 6'b001100;
frog_bram[324] = 6'b001100;
frog_bram[325] = 6'b000000;
frog_bram[326] = 6'b000000;
frog_bram[327] = 6'b000000;
frog_bram[328] = 6'b001100;
frog_bram[329] = 6'b001100;
frog_bram[330] = 6'b001100;
frog_bram[331] = 6'b001000;
frog_bram[332] = 6'b001000;
frog_bram[333] = 6'b001000;
frog_bram[334] = 6'b001100;
frog_bram[335] = 6'b001100;
frog_bram[336] = 6'b001100;
frog_bram[337] = 6'b001100;
frog_bram[338] = 6'b001100;
frog_bram[339] = 6'b001100;
frog_bram[340] = 6'b001100;
frog_bram[341] = 6'b001100;
frog_bram[342] = 6'b001100;
frog_bram[343] = 6'b001100;
frog_bram[344] = 6'b000000;
frog_bram[345] = 6'b000000;
frog_bram[346] = 6'b000000;
frog_bram[347] = 6'b001100;
frog_bram[348] = 6'b001100;
frog_bram[349] = 6'b001100;
frog_bram[350] = 6'b000000;
frog_bram[351] = 6'b000000;
frog_bram[352] = 6'b000000;
frog_bram[353] = 6'b000000;
frog_bram[354] = 6'b001100;
frog_bram[355] = 6'b001100;
frog_bram[356] = 6'b001100;
frog_bram[357] = 6'b001000;
frog_bram[358] = 6'b000000;
frog_bram[359] = 6'b000000;
frog_bram[360] = 6'b000000;
frog_bram[361] = 6'b001100;
frog_bram[362] = 6'b001100;
frog_bram[363] = 6'b001100;
frog_bram[364] = 6'b001100;
frog_bram[365] = 6'b001100;
frog_bram[366] = 6'b001100;
frog_bram[367] = 6'b001100;
frog_bram[368] = 6'b001100;
frog_bram[369] = 6'b001100;
frog_bram[370] = 6'b001100;
frog_bram[371] = 6'b001100;
frog_bram[372] = 6'b001100;
frog_bram[373] = 6'b001100;
frog_bram[374] = 6'b001100;
frog_bram[375] = 6'b000000;
frog_bram[376] = 6'b000000;
frog_bram[377] = 6'b000000;
frog_bram[378] = 6'b001000;
frog_bram[379] = 6'b001100;
frog_bram[380] = 6'b001100;
frog_bram[381] = 6'b001100;
frog_bram[382] = 6'b000000;
frog_bram[383] = 6'b000000;
frog_bram[384] = 6'b000000;
frog_bram[385] = 6'b000000;
frog_bram[386] = 6'b001100;
frog_bram[387] = 6'b001100;
frog_bram[388] = 6'b001100;
frog_bram[389] = 6'b001000;
frog_bram[390] = 6'b001000;
frog_bram[391] = 6'b001000;
frog_bram[392] = 6'b000000;
frog_bram[393] = 6'b000000;
frog_bram[394] = 6'b001000;
frog_bram[395] = 6'b001100;
frog_bram[396] = 6'b001100;
frog_bram[397] = 6'b001100;
frog_bram[398] = 6'b001100;
frog_bram[399] = 6'b001100;
frog_bram[400] = 6'b001100;
frog_bram[401] = 6'b001100;
frog_bram[402] = 6'b001100;
frog_bram[403] = 6'b001100;
frog_bram[404] = 6'b001100;
frog_bram[405] = 6'b001000;
frog_bram[406] = 6'b000000;
frog_bram[407] = 6'b000000;
frog_bram[408] = 6'b001000;
frog_bram[409] = 6'b001000;
frog_bram[410] = 6'b001000;
frog_bram[411] = 6'b001100;
frog_bram[412] = 6'b001100;
frog_bram[413] = 6'b001100;
frog_bram[414] = 6'b000000;
frog_bram[415] = 6'b000000;
frog_bram[416] = 6'b000000;
frog_bram[417] = 6'b000000;
frog_bram[418] = 6'b000000;
frog_bram[419] = 6'b001000;
frog_bram[420] = 6'b001000;
frog_bram[421] = 6'b001000;
frog_bram[422] = 6'b001000;
frog_bram[423] = 6'b001000;
frog_bram[424] = 6'b001000;
frog_bram[425] = 6'b000000;
frog_bram[426] = 6'b001000;
frog_bram[427] = 6'b001100;
frog_bram[428] = 6'b001100;
frog_bram[429] = 6'b001100;
frog_bram[430] = 6'b001000;
frog_bram[431] = 6'b001000;
frog_bram[432] = 6'b001000;
frog_bram[433] = 6'b001000;
frog_bram[434] = 6'b001100;
frog_bram[435] = 6'b001100;
frog_bram[436] = 6'b001100;
frog_bram[437] = 6'b001000;
frog_bram[438] = 6'b000000;
frog_bram[439] = 6'b001000;
frog_bram[440] = 6'b001000;
frog_bram[441] = 6'b001000;
frog_bram[442] = 6'b001000;
frog_bram[443] = 6'b001000;
frog_bram[444] = 6'b001000;
frog_bram[445] = 6'b000000;
frog_bram[446] = 6'b000000;
frog_bram[447] = 6'b000000;
frog_bram[448] = 6'b000000;
frog_bram[449] = 6'b000000;
frog_bram[450] = 6'b000000;
frog_bram[451] = 6'b000000;
frog_bram[452] = 6'b001000;
frog_bram[453] = 6'b001000;
frog_bram[454] = 6'b001000;
frog_bram[455] = 6'b001000;
frog_bram[456] = 6'b001100;
frog_bram[457] = 6'b001000;
frog_bram[458] = 6'b001100;
frog_bram[459] = 6'b001100;
frog_bram[460] = 6'b001100;
frog_bram[461] = 6'b001100;
frog_bram[462] = 6'b001100;
frog_bram[463] = 6'b001000;
frog_bram[464] = 6'b001000;
frog_bram[465] = 6'b001100;
frog_bram[466] = 6'b001100;
frog_bram[467] = 6'b001100;
frog_bram[468] = 6'b001100;
frog_bram[469] = 6'b001100;
frog_bram[470] = 6'b001000;
frog_bram[471] = 6'b001100;
frog_bram[472] = 6'b001000;
frog_bram[473] = 6'b001000;
frog_bram[474] = 6'b001000;
frog_bram[475] = 6'b001000;
frog_bram[476] = 6'b000000;
frog_bram[477] = 6'b000000;
frog_bram[478] = 6'b000000;
frog_bram[479] = 6'b000000;
frog_bram[480] = 6'b000000;
frog_bram[481] = 6'b000000;
frog_bram[482] = 6'b000000;
frog_bram[483] = 6'b000000;
frog_bram[484] = 6'b000000;
frog_bram[485] = 6'b000000;
frog_bram[486] = 6'b001000;
frog_bram[487] = 6'b001100;
frog_bram[488] = 6'b000000;
frog_bram[489] = 6'b001100;
frog_bram[490] = 6'b001100;
frog_bram[491] = 6'b001100;
frog_bram[492] = 6'b001100;
frog_bram[493] = 6'b001100;
frog_bram[494] = 6'b001100;
frog_bram[495] = 6'b001000;
frog_bram[496] = 6'b001000;
frog_bram[497] = 6'b001100;
frog_bram[498] = 6'b001100;
frog_bram[499] = 6'b001100;
frog_bram[500] = 6'b001100;
frog_bram[501] = 6'b001100;
frog_bram[502] = 6'b001100;
frog_bram[503] = 6'b000000;
frog_bram[504] = 6'b001100;
frog_bram[505] = 6'b001000;
frog_bram[506] = 6'b000000;
frog_bram[507] = 6'b000000;
frog_bram[508] = 6'b000000;
frog_bram[509] = 6'b000000;
frog_bram[510] = 6'b000000;
frog_bram[511] = 6'b000000;
frog_bram[512] = 6'b000000;
frog_bram[513] = 6'b000000;
frog_bram[514] = 6'b000000;
frog_bram[515] = 6'b000000;
frog_bram[516] = 6'b000000;
frog_bram[517] = 6'b000000;
frog_bram[518] = 6'b000000;
frog_bram[519] = 6'b001000;
frog_bram[520] = 6'b000000;
frog_bram[521] = 6'b001100;
frog_bram[522] = 6'b001100;
frog_bram[523] = 6'b001100;
frog_bram[524] = 6'b001100;
frog_bram[525] = 6'b001100;
frog_bram[526] = 6'b001000;
frog_bram[527] = 6'b001000;
frog_bram[528] = 6'b001000;
frog_bram[529] = 6'b001000;
frog_bram[530] = 6'b001100;
frog_bram[531] = 6'b001100;
frog_bram[532] = 6'b001100;
frog_bram[533] = 6'b001100;
frog_bram[534] = 6'b001100;
frog_bram[535] = 6'b000000;
frog_bram[536] = 6'b001000;
frog_bram[537] = 6'b000000;
frog_bram[538] = 6'b000000;
frog_bram[539] = 6'b000000;
frog_bram[540] = 6'b000000;
frog_bram[541] = 6'b000000;
frog_bram[542] = 6'b000000;
frog_bram[543] = 6'b000000;
frog_bram[544] = 6'b000000;
frog_bram[545] = 6'b000000;
frog_bram[546] = 6'b000000;
frog_bram[547] = 6'b000000;
frog_bram[548] = 6'b000000;
frog_bram[549] = 6'b000000;
frog_bram[550] = 6'b000000;
frog_bram[551] = 6'b000000;
frog_bram[552] = 6'b001000;
frog_bram[553] = 6'b001100;
frog_bram[554] = 6'b001100;
frog_bram[555] = 6'b001100;
frog_bram[556] = 6'b001100;
frog_bram[557] = 6'b001000;
frog_bram[558] = 6'b001000;
frog_bram[559] = 6'b001000;
frog_bram[560] = 6'b001000;
frog_bram[561] = 6'b001000;
frog_bram[562] = 6'b001000;
frog_bram[563] = 6'b001100;
frog_bram[564] = 6'b001100;
frog_bram[565] = 6'b001100;
frog_bram[566] = 6'b001100;
frog_bram[567] = 6'b001000;
frog_bram[568] = 6'b000000;
frog_bram[569] = 6'b000000;
frog_bram[570] = 6'b000000;
frog_bram[571] = 6'b000000;
frog_bram[572] = 6'b000000;
frog_bram[573] = 6'b000000;
frog_bram[574] = 6'b000000;
frog_bram[575] = 6'b000000;
frog_bram[576] = 6'b000000;
frog_bram[577] = 6'b000000;
frog_bram[578] = 6'b000000;
frog_bram[579] = 6'b000000;
frog_bram[580] = 6'b000000;
frog_bram[581] = 6'b000000;
frog_bram[582] = 6'b001000;
frog_bram[583] = 6'b001000;
frog_bram[584] = 6'b000000;
frog_bram[585] = 6'b001100;
frog_bram[586] = 6'b001100;
frog_bram[587] = 6'b001100;
frog_bram[588] = 6'b001100;
frog_bram[589] = 6'b001100;
frog_bram[590] = 6'b001000;
frog_bram[591] = 6'b001000;
frog_bram[592] = 6'b001000;
frog_bram[593] = 6'b001000;
frog_bram[594] = 6'b001100;
frog_bram[595] = 6'b001100;
frog_bram[596] = 6'b001100;
frog_bram[597] = 6'b001100;
frog_bram[598] = 6'b001100;
frog_bram[599] = 6'b000000;
frog_bram[600] = 6'b001000;
frog_bram[601] = 6'b001000;
frog_bram[602] = 6'b000000;
frog_bram[603] = 6'b000000;
frog_bram[604] = 6'b000000;
frog_bram[605] = 6'b000000;
frog_bram[606] = 6'b000000;
frog_bram[607] = 6'b000000;
frog_bram[608] = 6'b000000;
frog_bram[609] = 6'b000000;
frog_bram[610] = 6'b000000;
frog_bram[611] = 6'b000000;
frog_bram[612] = 6'b000000;
frog_bram[613] = 6'b001000;
frog_bram[614] = 6'b001100;
frog_bram[615] = 6'b001000;
frog_bram[616] = 6'b000000;
frog_bram[617] = 6'b001100;
frog_bram[618] = 6'b001100;
frog_bram[619] = 6'b001100;
frog_bram[620] = 6'b001100;
frog_bram[621] = 6'b001100;
frog_bram[622] = 6'b001000;
frog_bram[623] = 6'b001000;
frog_bram[624] = 6'b001000;
frog_bram[625] = 6'b001000;
frog_bram[626] = 6'b001100;
frog_bram[627] = 6'b001100;
frog_bram[628] = 6'b001100;
frog_bram[629] = 6'b001100;
frog_bram[630] = 6'b001100;
frog_bram[631] = 6'b000000;
frog_bram[632] = 6'b001000;
frog_bram[633] = 6'b001100;
frog_bram[634] = 6'b001000;
frog_bram[635] = 6'b000000;
frog_bram[636] = 6'b000000;
frog_bram[637] = 6'b000000;
frog_bram[638] = 6'b000000;
frog_bram[639] = 6'b000000;
frog_bram[640] = 6'b000000;
frog_bram[641] = 6'b000000;
frog_bram[642] = 6'b000000;
frog_bram[643] = 6'b000000;
frog_bram[644] = 6'b000000;
frog_bram[645] = 6'b001000;
frog_bram[646] = 6'b001100;
frog_bram[647] = 6'b001000;
frog_bram[648] = 6'b000000;
frog_bram[649] = 6'b001000;
frog_bram[650] = 6'b001100;
frog_bram[651] = 6'b001100;
frog_bram[652] = 6'b001100;
frog_bram[653] = 6'b001100;
frog_bram[654] = 6'b001000;
frog_bram[655] = 6'b001000;
frog_bram[656] = 6'b001000;
frog_bram[657] = 6'b001000;
frog_bram[658] = 6'b001100;
frog_bram[659] = 6'b001100;
frog_bram[660] = 6'b001100;
frog_bram[661] = 6'b001100;
frog_bram[662] = 6'b001000;
frog_bram[663] = 6'b000000;
frog_bram[664] = 6'b001000;
frog_bram[665] = 6'b001100;
frog_bram[666] = 6'b001000;
frog_bram[667] = 6'b000000;
frog_bram[668] = 6'b000000;
frog_bram[669] = 6'b000000;
frog_bram[670] = 6'b000000;
frog_bram[671] = 6'b000000;
frog_bram[672] = 6'b000000;
frog_bram[673] = 6'b000000;
frog_bram[674] = 6'b000000;
frog_bram[675] = 6'b000000;
frog_bram[676] = 6'b000000;
frog_bram[677] = 6'b001000;
frog_bram[678] = 6'b001100;
frog_bram[679] = 6'b001000;
frog_bram[680] = 6'b000000;
frog_bram[681] = 6'b001000;
frog_bram[682] = 6'b001100;
frog_bram[683] = 6'b001100;
frog_bram[684] = 6'b001000;
frog_bram[685] = 6'b001000;
frog_bram[686] = 6'b001000;
frog_bram[687] = 6'b001000;
frog_bram[688] = 6'b001000;
frog_bram[689] = 6'b001000;
frog_bram[690] = 6'b001000;
frog_bram[691] = 6'b001000;
frog_bram[692] = 6'b001100;
frog_bram[693] = 6'b001100;
frog_bram[694] = 6'b001000;
frog_bram[695] = 6'b000000;
frog_bram[696] = 6'b001000;
frog_bram[697] = 6'b001100;
frog_bram[698] = 6'b001000;
frog_bram[699] = 6'b000000;
frog_bram[700] = 6'b000000;
frog_bram[701] = 6'b000000;
frog_bram[702] = 6'b000000;
frog_bram[703] = 6'b000000;
frog_bram[704] = 6'b000000;
frog_bram[705] = 6'b000000;
frog_bram[706] = 6'b001000;
frog_bram[707] = 6'b001000;
frog_bram[708] = 6'b000000;
frog_bram[709] = 6'b001000;
frog_bram[710] = 6'b001100;
frog_bram[711] = 6'b001100;
frog_bram[712] = 6'b001000;
frog_bram[713] = 6'b000000;
frog_bram[714] = 6'b001000;
frog_bram[715] = 6'b001000;
frog_bram[716] = 6'b001000;
frog_bram[717] = 6'b001000;
frog_bram[718] = 6'b001000;
frog_bram[719] = 6'b001000;
frog_bram[720] = 6'b001000;
frog_bram[721] = 6'b001000;
frog_bram[722] = 6'b001000;
frog_bram[723] = 6'b001000;
frog_bram[724] = 6'b001000;
frog_bram[725] = 6'b001000;
frog_bram[726] = 6'b000000;
frog_bram[727] = 6'b001000;
frog_bram[728] = 6'b001100;
frog_bram[729] = 6'b001100;
frog_bram[730] = 6'b001000;
frog_bram[731] = 6'b000000;
frog_bram[732] = 6'b001000;
frog_bram[733] = 6'b001000;
frog_bram[734] = 6'b000000;
frog_bram[735] = 6'b000000;
frog_bram[736] = 6'b000000;
frog_bram[737] = 6'b000000;
frog_bram[738] = 6'b001100;
frog_bram[739] = 6'b001100;
frog_bram[740] = 6'b000000;
frog_bram[741] = 6'b001000;
frog_bram[742] = 6'b001100;
frog_bram[743] = 6'b001100;
frog_bram[744] = 6'b001000;
frog_bram[745] = 6'b000000;
frog_bram[746] = 6'b001000;
frog_bram[747] = 6'b001100;
frog_bram[748] = 6'b001100;
frog_bram[749] = 6'b001100;
frog_bram[750] = 6'b001000;
frog_bram[751] = 6'b001000;
frog_bram[752] = 6'b001000;
frog_bram[753] = 6'b001000;
frog_bram[754] = 6'b001100;
frog_bram[755] = 6'b001100;
frog_bram[756] = 6'b001100;
frog_bram[757] = 6'b001000;
frog_bram[758] = 6'b000000;
frog_bram[759] = 6'b001000;
frog_bram[760] = 6'b001100;
frog_bram[761] = 6'b001100;
frog_bram[762] = 6'b001000;
frog_bram[763] = 6'b000000;
frog_bram[764] = 6'b001100;
frog_bram[765] = 6'b001100;
frog_bram[766] = 6'b000000;
frog_bram[767] = 6'b000000;
frog_bram[768] = 6'b001000;
frog_bram[769] = 6'b001000;
frog_bram[770] = 6'b000100;
frog_bram[771] = 6'b001100;
frog_bram[772] = 6'b000000;
frog_bram[773] = 6'b001000;
frog_bram[774] = 6'b001000;
frog_bram[775] = 6'b001100;
frog_bram[776] = 6'b001000;
frog_bram[777] = 6'b000000;
frog_bram[778] = 6'b001000;
frog_bram[779] = 6'b001100;
frog_bram[780] = 6'b001100;
frog_bram[781] = 6'b001100;
frog_bram[782] = 6'b001000;
frog_bram[783] = 6'b001000;
frog_bram[784] = 6'b001000;
frog_bram[785] = 6'b001000;
frog_bram[786] = 6'b001100;
frog_bram[787] = 6'b001100;
frog_bram[788] = 6'b001100;
frog_bram[789] = 6'b001000;
frog_bram[790] = 6'b000000;
frog_bram[791] = 6'b001000;
frog_bram[792] = 6'b001100;
frog_bram[793] = 6'b001000;
frog_bram[794] = 6'b001000;
frog_bram[795] = 6'b000000;
frog_bram[796] = 6'b001100;
frog_bram[797] = 6'b000100;
frog_bram[798] = 6'b001000;
frog_bram[799] = 6'b001000;
frog_bram[800] = 6'b001100;
frog_bram[801] = 6'b001100;
frog_bram[802] = 6'b001000;
frog_bram[803] = 6'b001100;
frog_bram[804] = 6'b001000;
frog_bram[805] = 6'b000000;
frog_bram[806] = 6'b001000;
frog_bram[807] = 6'b001100;
frog_bram[808] = 6'b001100;
frog_bram[809] = 6'b001000;
frog_bram[810] = 6'b000000;
frog_bram[811] = 6'b001000;
frog_bram[812] = 6'b001100;
frog_bram[813] = 6'b001000;
frog_bram[814] = 6'b001000;
frog_bram[815] = 6'b001000;
frog_bram[816] = 6'b001000;
frog_bram[817] = 6'b001000;
frog_bram[818] = 6'b001000;
frog_bram[819] = 6'b001100;
frog_bram[820] = 6'b001000;
frog_bram[821] = 6'b000000;
frog_bram[822] = 6'b001000;
frog_bram[823] = 6'b001100;
frog_bram[824] = 6'b001100;
frog_bram[825] = 6'b001000;
frog_bram[826] = 6'b000000;
frog_bram[827] = 6'b001000;
frog_bram[828] = 6'b001100;
frog_bram[829] = 6'b001000;
frog_bram[830] = 6'b001100;
frog_bram[831] = 6'b001100;
frog_bram[832] = 6'b000000;
frog_bram[833] = 6'b001100;
frog_bram[834] = 6'b001100;
frog_bram[835] = 6'b001100;
frog_bram[836] = 6'b001100;
frog_bram[837] = 6'b001000;
frog_bram[838] = 6'b000000;
frog_bram[839] = 6'b001100;
frog_bram[840] = 6'b001100;
frog_bram[841] = 6'b001000;
frog_bram[842] = 6'b000000;
frog_bram[843] = 6'b001000;
frog_bram[844] = 6'b001000;
frog_bram[845] = 6'b001000;
frog_bram[846] = 6'b001000;
frog_bram[847] = 6'b001000;
frog_bram[848] = 6'b001000;
frog_bram[849] = 6'b001000;
frog_bram[850] = 6'b001000;
frog_bram[851] = 6'b001000;
frog_bram[852] = 6'b001000;
frog_bram[853] = 6'b000000;
frog_bram[854] = 6'b001000;
frog_bram[855] = 6'b001100;
frog_bram[856] = 6'b001100;
frog_bram[857] = 6'b000000;
frog_bram[858] = 6'b001000;
frog_bram[859] = 6'b001100;
frog_bram[860] = 6'b001100;
frog_bram[861] = 6'b001100;
frog_bram[862] = 6'b001100;
frog_bram[863] = 6'b000000;
frog_bram[864] = 6'b001000;
frog_bram[865] = 6'b001100;
frog_bram[866] = 6'b001100;
frog_bram[867] = 6'b001100;
frog_bram[868] = 6'b001100;
frog_bram[869] = 6'b001100;
frog_bram[870] = 6'b001100;
frog_bram[871] = 6'b001100;
frog_bram[872] = 6'b001100;
frog_bram[873] = 6'b001000;
frog_bram[874] = 6'b000000;
frog_bram[875] = 6'b000000;
frog_bram[876] = 6'b000000;
frog_bram[877] = 6'b001000;
frog_bram[878] = 6'b001000;
frog_bram[879] = 6'b001000;
frog_bram[880] = 6'b001000;
frog_bram[881] = 6'b001000;
frog_bram[882] = 6'b001000;
frog_bram[883] = 6'b000000;
frog_bram[884] = 6'b000000;
frog_bram[885] = 6'b000000;
frog_bram[886] = 6'b001000;
frog_bram[887] = 6'b001100;
frog_bram[888] = 6'b001100;
frog_bram[889] = 6'b001100;
frog_bram[890] = 6'b001100;
frog_bram[891] = 6'b001100;
frog_bram[892] = 6'b001100;
frog_bram[893] = 6'b001100;
frog_bram[894] = 6'b001100;
frog_bram[895] = 6'b001000;
frog_bram[896] = 6'b001100;
frog_bram[897] = 6'b001100;
frog_bram[898] = 6'b001100;
frog_bram[899] = 6'b001100;
frog_bram[900] = 6'b001100;
frog_bram[901] = 6'b001100;
frog_bram[902] = 6'b001100;
frog_bram[903] = 6'b001100;
frog_bram[904] = 6'b001100;
frog_bram[905] = 6'b000000;
frog_bram[906] = 6'b000000;
frog_bram[907] = 6'b000000;
frog_bram[908] = 6'b000000;
frog_bram[909] = 6'b000000;
frog_bram[910] = 6'b000000;
frog_bram[911] = 6'b001000;
frog_bram[912] = 6'b001000;
frog_bram[913] = 6'b000000;
frog_bram[914] = 6'b000000;
frog_bram[915] = 6'b000000;
frog_bram[916] = 6'b000000;
frog_bram[917] = 6'b000000;
frog_bram[918] = 6'b000000;
frog_bram[919] = 6'b001100;
frog_bram[920] = 6'b001100;
frog_bram[921] = 6'b001100;
frog_bram[922] = 6'b001100;
frog_bram[923] = 6'b001100;
frog_bram[924] = 6'b001100;
frog_bram[925] = 6'b001100;
frog_bram[926] = 6'b001100;
frog_bram[927] = 6'b001100;
frog_bram[928] = 6'b000000;
frog_bram[929] = 6'b000000;
frog_bram[930] = 6'b001000;
frog_bram[931] = 6'b001000;
frog_bram[932] = 6'b001000;
frog_bram[933] = 6'b001100;
frog_bram[934] = 6'b001100;
frog_bram[935] = 6'b001100;
frog_bram[936] = 6'b001000;
frog_bram[937] = 6'b000000;
frog_bram[938] = 6'b000000;
frog_bram[939] = 6'b000000;
frog_bram[940] = 6'b000000;
frog_bram[941] = 6'b000000;
frog_bram[942] = 6'b000000;
frog_bram[943] = 6'b000000;
frog_bram[944] = 6'b000000;
frog_bram[945] = 6'b000000;
frog_bram[946] = 6'b000000;
frog_bram[947] = 6'b000000;
frog_bram[948] = 6'b000000;
frog_bram[949] = 6'b000000;
frog_bram[950] = 6'b000000;
frog_bram[951] = 6'b001000;
frog_bram[952] = 6'b001100;
frog_bram[953] = 6'b001100;
frog_bram[954] = 6'b001100;
frog_bram[955] = 6'b001000;
frog_bram[956] = 6'b001000;
frog_bram[957] = 6'b001000;
frog_bram[958] = 6'b000000;
frog_bram[959] = 6'b000000;
frog_bram[960] = 6'b000000;
frog_bram[961] = 6'b000000;
frog_bram[962] = 6'b000000;
frog_bram[963] = 6'b000000;
frog_bram[964] = 6'b000000;
frog_bram[965] = 6'b001000;
frog_bram[966] = 6'b001000;
frog_bram[967] = 6'b000000;
frog_bram[968] = 6'b000000;
frog_bram[969] = 6'b000000;
frog_bram[970] = 6'b000000;
frog_bram[971] = 6'b000000;
frog_bram[972] = 6'b000000;
frog_bram[973] = 6'b000000;
frog_bram[974] = 6'b000000;
frog_bram[975] = 6'b000000;
frog_bram[976] = 6'b000000;
frog_bram[977] = 6'b000000;
frog_bram[978] = 6'b000000;
frog_bram[979] = 6'b000000;
frog_bram[980] = 6'b000000;
frog_bram[981] = 6'b000000;
frog_bram[982] = 6'b000000;
frog_bram[983] = 6'b000000;
frog_bram[984] = 6'b000000;
frog_bram[985] = 6'b001000;
frog_bram[986] = 6'b001000;
frog_bram[987] = 6'b000000;
frog_bram[988] = 6'b000000;
frog_bram[989] = 6'b000000;
frog_bram[990] = 6'b000000;
frog_bram[991] = 6'b000000;
frog_bram[992] = 6'b000000;
frog_bram[993] = 6'b000000;
frog_bram[994] = 6'b000000;
frog_bram[995] = 6'b000000;
frog_bram[996] = 6'b000000;
frog_bram[997] = 6'b000000;
frog_bram[998] = 6'b000000;
frog_bram[999] = 6'b000000;
frog_bram[1000] = 6'b000000;
frog_bram[1001] = 6'b000000;
frog_bram[1002] = 6'b000000;
frog_bram[1003] = 6'b000000;
frog_bram[1004] = 6'b000000;
frog_bram[1005] = 6'b000000;
frog_bram[1006] = 6'b000000;
frog_bram[1007] = 6'b000000;
frog_bram[1008] = 6'b000000;
frog_bram[1009] = 6'b000000;
frog_bram[1010] = 6'b000000;
frog_bram[1011] = 6'b000000;
frog_bram[1012] = 6'b000000;
frog_bram[1013] = 6'b000000;
frog_bram[1014] = 6'b000000;
frog_bram[1015] = 6'b000000;
frog_bram[1016] = 6'b000000;
frog_bram[1017] = 6'b000000;
frog_bram[1018] = 6'b000000;
frog_bram[1019] = 6'b000000;
frog_bram[1020] = 6'b000000;
frog_bram[1021] = 6'b000000;
frog_bram[1022] = 6'b000000;
frog_bram[1023] = 6'b000000;
        // Add more initialization here for the down-facing sprite (1024 - 2047)
frog_bram[1024] = 6'b000000;
frog_bram[1025] = 6'b000000;
frog_bram[1026] = 6'b000000;
frog_bram[1027] = 6'b000000;
frog_bram[1028] = 6'b000000;
frog_bram[1029] = 6'b000000;
frog_bram[1030] = 6'b000000;
frog_bram[1031] = 6'b000000;
frog_bram[1032] = 6'b000000;
frog_bram[1033] = 6'b000000;
frog_bram[1034] = 6'b000000;
frog_bram[1035] = 6'b000000;
frog_bram[1036] = 6'b000000;
frog_bram[1037] = 6'b000000;
frog_bram[1038] = 6'b000000;
frog_bram[1039] = 6'b000000;
frog_bram[1040] = 6'b000000;
frog_bram[1041] = 6'b000000;
frog_bram[1042] = 6'b000000;
frog_bram[1043] = 6'b000000;
frog_bram[1044] = 6'b000000;
frog_bram[1045] = 6'b000000;
frog_bram[1046] = 6'b000000;
frog_bram[1047] = 6'b000000;
frog_bram[1048] = 6'b000000;
frog_bram[1049] = 6'b000000;
frog_bram[1050] = 6'b000000;
frog_bram[1051] = 6'b000000;
frog_bram[1052] = 6'b000000;
frog_bram[1053] = 6'b000000;
frog_bram[1054] = 6'b000000;
frog_bram[1055] = 6'b000000;
frog_bram[1056] = 6'b000000;
frog_bram[1057] = 6'b000000;
frog_bram[1058] = 6'b000000;
frog_bram[1059] = 6'b000000;
frog_bram[1060] = 6'b000000;
frog_bram[1061] = 6'b001000;
frog_bram[1062] = 6'b001000;
frog_bram[1063] = 6'b000000;
frog_bram[1064] = 6'b000000;
frog_bram[1065] = 6'b000000;
frog_bram[1066] = 6'b000000;
frog_bram[1067] = 6'b000000;
frog_bram[1068] = 6'b000000;
frog_bram[1069] = 6'b000000;
frog_bram[1070] = 6'b000000;
frog_bram[1071] = 6'b000000;
frog_bram[1072] = 6'b000000;
frog_bram[1073] = 6'b000000;
frog_bram[1074] = 6'b000000;
frog_bram[1075] = 6'b000000;
frog_bram[1076] = 6'b000000;
frog_bram[1077] = 6'b000000;
frog_bram[1078] = 6'b000000;
frog_bram[1079] = 6'b000000;
frog_bram[1080] = 6'b000000;
frog_bram[1081] = 6'b001000;
frog_bram[1082] = 6'b001000;
frog_bram[1083] = 6'b000000;
frog_bram[1084] = 6'b000000;
frog_bram[1085] = 6'b000000;
frog_bram[1086] = 6'b000000;
frog_bram[1087] = 6'b000000;
frog_bram[1088] = 6'b000000;
frog_bram[1089] = 6'b000000;
frog_bram[1090] = 6'b001000;
frog_bram[1091] = 6'b001000;
frog_bram[1092] = 6'b001000;
frog_bram[1093] = 6'b001100;
frog_bram[1094] = 6'b001100;
frog_bram[1095] = 6'b001100;
frog_bram[1096] = 6'b001000;
frog_bram[1097] = 6'b000000;
frog_bram[1098] = 6'b000000;
frog_bram[1099] = 6'b000000;
frog_bram[1100] = 6'b000000;
frog_bram[1101] = 6'b000000;
frog_bram[1102] = 6'b000000;
frog_bram[1103] = 6'b000000;
frog_bram[1104] = 6'b000000;
frog_bram[1105] = 6'b000000;
frog_bram[1106] = 6'b000000;
frog_bram[1107] = 6'b000000;
frog_bram[1108] = 6'b000000;
frog_bram[1109] = 6'b000000;
frog_bram[1110] = 6'b000000;
frog_bram[1111] = 6'b001000;
frog_bram[1112] = 6'b001100;
frog_bram[1113] = 6'b001100;
frog_bram[1114] = 6'b001100;
frog_bram[1115] = 6'b001000;
frog_bram[1116] = 6'b001000;
frog_bram[1117] = 6'b001000;
frog_bram[1118] = 6'b000000;
frog_bram[1119] = 6'b000000;
frog_bram[1120] = 6'b001100;
frog_bram[1121] = 6'b001100;
frog_bram[1122] = 6'b001100;
frog_bram[1123] = 6'b001100;
frog_bram[1124] = 6'b001100;
frog_bram[1125] = 6'b001100;
frog_bram[1126] = 6'b001100;
frog_bram[1127] = 6'b001100;
frog_bram[1128] = 6'b001100;
frog_bram[1129] = 6'b000000;
frog_bram[1130] = 6'b000000;
frog_bram[1131] = 6'b000000;
frog_bram[1132] = 6'b000000;
frog_bram[1133] = 6'b000000;
frog_bram[1134] = 6'b000000;
frog_bram[1135] = 6'b001000;
frog_bram[1136] = 6'b001000;
frog_bram[1137] = 6'b000000;
frog_bram[1138] = 6'b000000;
frog_bram[1139] = 6'b000000;
frog_bram[1140] = 6'b000000;
frog_bram[1141] = 6'b000000;
frog_bram[1142] = 6'b000000;
frog_bram[1143] = 6'b001100;
frog_bram[1144] = 6'b001100;
frog_bram[1145] = 6'b001100;
frog_bram[1146] = 6'b001100;
frog_bram[1147] = 6'b001100;
frog_bram[1148] = 6'b001100;
frog_bram[1149] = 6'b001100;
frog_bram[1150] = 6'b001100;
frog_bram[1151] = 6'b001100;
frog_bram[1152] = 6'b001000;
frog_bram[1153] = 6'b001100;
frog_bram[1154] = 6'b001100;
frog_bram[1155] = 6'b001100;
frog_bram[1156] = 6'b001100;
frog_bram[1157] = 6'b001100;
frog_bram[1158] = 6'b001100;
frog_bram[1159] = 6'b001100;
frog_bram[1160] = 6'b001100;
frog_bram[1161] = 6'b001000;
frog_bram[1162] = 6'b000000;
frog_bram[1163] = 6'b000000;
frog_bram[1164] = 6'b000000;
frog_bram[1165] = 6'b001000;
frog_bram[1166] = 6'b001000;
frog_bram[1167] = 6'b001000;
frog_bram[1168] = 6'b001000;
frog_bram[1169] = 6'b001000;
frog_bram[1170] = 6'b001000;
frog_bram[1171] = 6'b000000;
frog_bram[1172] = 6'b000000;
frog_bram[1173] = 6'b000000;
frog_bram[1174] = 6'b001000;
frog_bram[1175] = 6'b001100;
frog_bram[1176] = 6'b001100;
frog_bram[1177] = 6'b001100;
frog_bram[1178] = 6'b001100;
frog_bram[1179] = 6'b001100;
frog_bram[1180] = 6'b001100;
frog_bram[1181] = 6'b001100;
frog_bram[1182] = 6'b001100;
frog_bram[1183] = 6'b001000;
frog_bram[1184] = 6'b000000;
frog_bram[1185] = 6'b001100;
frog_bram[1186] = 6'b001100;
frog_bram[1187] = 6'b001100;
frog_bram[1188] = 6'b001100;
frog_bram[1189] = 6'b001000;
frog_bram[1190] = 6'b000000;
frog_bram[1191] = 6'b001100;
frog_bram[1192] = 6'b001100;
frog_bram[1193] = 6'b001000;
frog_bram[1194] = 6'b000000;
frog_bram[1195] = 6'b001000;
frog_bram[1196] = 6'b001000;
frog_bram[1197] = 6'b001000;
frog_bram[1198] = 6'b001000;
frog_bram[1199] = 6'b001000;
frog_bram[1200] = 6'b001000;
frog_bram[1201] = 6'b001000;
frog_bram[1202] = 6'b001000;
frog_bram[1203] = 6'b001000;
frog_bram[1204] = 6'b001000;
frog_bram[1205] = 6'b000000;
frog_bram[1206] = 6'b001000;
frog_bram[1207] = 6'b001100;
frog_bram[1208] = 6'b001100;
frog_bram[1209] = 6'b000000;
frog_bram[1210] = 6'b001000;
frog_bram[1211] = 6'b001100;
frog_bram[1212] = 6'b001100;
frog_bram[1213] = 6'b001100;
frog_bram[1214] = 6'b001100;
frog_bram[1215] = 6'b000000;
frog_bram[1216] = 6'b001100;
frog_bram[1217] = 6'b001100;
frog_bram[1218] = 6'b001000;
frog_bram[1219] = 6'b001100;
frog_bram[1220] = 6'b001000;
frog_bram[1221] = 6'b000000;
frog_bram[1222] = 6'b001000;
frog_bram[1223] = 6'b001100;
frog_bram[1224] = 6'b001100;
frog_bram[1225] = 6'b001000;
frog_bram[1226] = 6'b000000;
frog_bram[1227] = 6'b001000;
frog_bram[1228] = 6'b001100;
frog_bram[1229] = 6'b001000;
frog_bram[1230] = 6'b001000;
frog_bram[1231] = 6'b001000;
frog_bram[1232] = 6'b001000;
frog_bram[1233] = 6'b001000;
frog_bram[1234] = 6'b001000;
frog_bram[1235] = 6'b001100;
frog_bram[1236] = 6'b001000;
frog_bram[1237] = 6'b000000;
frog_bram[1238] = 6'b001000;
frog_bram[1239] = 6'b001100;
frog_bram[1240] = 6'b001100;
frog_bram[1241] = 6'b001000;
frog_bram[1242] = 6'b000000;
frog_bram[1243] = 6'b001000;
frog_bram[1244] = 6'b001100;
frog_bram[1245] = 6'b001000;
frog_bram[1246] = 6'b001100;
frog_bram[1247] = 6'b001100;
frog_bram[1248] = 6'b001000;
frog_bram[1249] = 6'b001000;
frog_bram[1250] = 6'b000100;
frog_bram[1251] = 6'b001100;
frog_bram[1252] = 6'b000000;
frog_bram[1253] = 6'b001000;
frog_bram[1254] = 6'b001000;
frog_bram[1255] = 6'b001100;
frog_bram[1256] = 6'b001000;
frog_bram[1257] = 6'b000000;
frog_bram[1258] = 6'b001000;
frog_bram[1259] = 6'b001100;
frog_bram[1260] = 6'b001100;
frog_bram[1261] = 6'b001100;
frog_bram[1262] = 6'b001000;
frog_bram[1263] = 6'b001000;
frog_bram[1264] = 6'b001000;
frog_bram[1265] = 6'b001000;
frog_bram[1266] = 6'b001100;
frog_bram[1267] = 6'b001100;
frog_bram[1268] = 6'b001100;
frog_bram[1269] = 6'b001000;
frog_bram[1270] = 6'b000000;
frog_bram[1271] = 6'b001000;
frog_bram[1272] = 6'b001100;
frog_bram[1273] = 6'b001000;
frog_bram[1274] = 6'b001000;
frog_bram[1275] = 6'b000000;
frog_bram[1276] = 6'b001100;
frog_bram[1277] = 6'b000100;
frog_bram[1278] = 6'b001000;
frog_bram[1279] = 6'b001000;
frog_bram[1280] = 6'b000000;
frog_bram[1281] = 6'b000000;
frog_bram[1282] = 6'b001100;
frog_bram[1283] = 6'b001100;
frog_bram[1284] = 6'b000000;
frog_bram[1285] = 6'b001000;
frog_bram[1286] = 6'b001100;
frog_bram[1287] = 6'b001100;
frog_bram[1288] = 6'b001000;
frog_bram[1289] = 6'b000000;
frog_bram[1290] = 6'b001000;
frog_bram[1291] = 6'b001100;
frog_bram[1292] = 6'b001100;
frog_bram[1293] = 6'b001100;
frog_bram[1294] = 6'b001000;
frog_bram[1295] = 6'b001000;
frog_bram[1296] = 6'b001000;
frog_bram[1297] = 6'b001000;
frog_bram[1298] = 6'b001100;
frog_bram[1299] = 6'b001100;
frog_bram[1300] = 6'b001100;
frog_bram[1301] = 6'b001000;
frog_bram[1302] = 6'b000000;
frog_bram[1303] = 6'b001000;
frog_bram[1304] = 6'b001100;
frog_bram[1305] = 6'b001100;
frog_bram[1306] = 6'b001000;
frog_bram[1307] = 6'b000000;
frog_bram[1308] = 6'b001100;
frog_bram[1309] = 6'b001100;
frog_bram[1310] = 6'b000000;
frog_bram[1311] = 6'b000000;
frog_bram[1312] = 6'b000000;
frog_bram[1313] = 6'b000000;
frog_bram[1314] = 6'b001000;
frog_bram[1315] = 6'b001000;
frog_bram[1316] = 6'b000000;
frog_bram[1317] = 6'b001000;
frog_bram[1318] = 6'b001100;
frog_bram[1319] = 6'b001100;
frog_bram[1320] = 6'b001000;
frog_bram[1321] = 6'b000000;
frog_bram[1322] = 6'b001000;
frog_bram[1323] = 6'b001000;
frog_bram[1324] = 6'b001000;
frog_bram[1325] = 6'b001000;
frog_bram[1326] = 6'b001000;
frog_bram[1327] = 6'b001000;
frog_bram[1328] = 6'b001000;
frog_bram[1329] = 6'b001000;
frog_bram[1330] = 6'b001000;
frog_bram[1331] = 6'b001000;
frog_bram[1332] = 6'b001000;
frog_bram[1333] = 6'b001000;
frog_bram[1334] = 6'b000000;
frog_bram[1335] = 6'b001000;
frog_bram[1336] = 6'b001100;
frog_bram[1337] = 6'b001100;
frog_bram[1338] = 6'b001000;
frog_bram[1339] = 6'b000000;
frog_bram[1340] = 6'b001000;
frog_bram[1341] = 6'b001000;
frog_bram[1342] = 6'b000000;
frog_bram[1343] = 6'b000000;
frog_bram[1344] = 6'b000000;
frog_bram[1345] = 6'b000000;
frog_bram[1346] = 6'b000000;
frog_bram[1347] = 6'b000000;
frog_bram[1348] = 6'b000000;
frog_bram[1349] = 6'b001000;
frog_bram[1350] = 6'b001100;
frog_bram[1351] = 6'b001000;
frog_bram[1352] = 6'b000000;
frog_bram[1353] = 6'b001000;
frog_bram[1354] = 6'b001100;
frog_bram[1355] = 6'b001100;
frog_bram[1356] = 6'b001000;
frog_bram[1357] = 6'b001000;
frog_bram[1358] = 6'b001000;
frog_bram[1359] = 6'b001000;
frog_bram[1360] = 6'b001000;
frog_bram[1361] = 6'b001000;
frog_bram[1362] = 6'b001000;
frog_bram[1363] = 6'b001000;
frog_bram[1364] = 6'b001100;
frog_bram[1365] = 6'b001100;
frog_bram[1366] = 6'b001000;
frog_bram[1367] = 6'b000000;
frog_bram[1368] = 6'b001000;
frog_bram[1369] = 6'b001100;
frog_bram[1370] = 6'b001000;
frog_bram[1371] = 6'b000000;
frog_bram[1372] = 6'b000000;
frog_bram[1373] = 6'b000000;
frog_bram[1374] = 6'b000000;
frog_bram[1375] = 6'b000000;
frog_bram[1376] = 6'b000000;
frog_bram[1377] = 6'b000000;
frog_bram[1378] = 6'b000000;
frog_bram[1379] = 6'b000000;
frog_bram[1380] = 6'b000000;
frog_bram[1381] = 6'b001000;
frog_bram[1382] = 6'b001100;
frog_bram[1383] = 6'b001000;
frog_bram[1384] = 6'b000000;
frog_bram[1385] = 6'b001000;
frog_bram[1386] = 6'b001100;
frog_bram[1387] = 6'b001100;
frog_bram[1388] = 6'b001100;
frog_bram[1389] = 6'b001100;
frog_bram[1390] = 6'b001000;
frog_bram[1391] = 6'b001000;
frog_bram[1392] = 6'b001000;
frog_bram[1393] = 6'b001000;
frog_bram[1394] = 6'b001100;
frog_bram[1395] = 6'b001100;
frog_bram[1396] = 6'b001100;
frog_bram[1397] = 6'b001100;
frog_bram[1398] = 6'b001000;
frog_bram[1399] = 6'b000000;
frog_bram[1400] = 6'b001000;
frog_bram[1401] = 6'b001100;
frog_bram[1402] = 6'b001000;
frog_bram[1403] = 6'b000000;
frog_bram[1404] = 6'b000000;
frog_bram[1405] = 6'b000000;
frog_bram[1406] = 6'b000000;
frog_bram[1407] = 6'b000000;
frog_bram[1408] = 6'b000000;
frog_bram[1409] = 6'b000000;
frog_bram[1410] = 6'b000000;
frog_bram[1411] = 6'b000000;
frog_bram[1412] = 6'b000000;
frog_bram[1413] = 6'b001000;
frog_bram[1414] = 6'b001100;
frog_bram[1415] = 6'b001000;
frog_bram[1416] = 6'b000000;
frog_bram[1417] = 6'b001100;
frog_bram[1418] = 6'b001100;
frog_bram[1419] = 6'b001100;
frog_bram[1420] = 6'b001100;
frog_bram[1421] = 6'b001100;
frog_bram[1422] = 6'b001000;
frog_bram[1423] = 6'b001000;
frog_bram[1424] = 6'b001000;
frog_bram[1425] = 6'b001000;
frog_bram[1426] = 6'b001100;
frog_bram[1427] = 6'b001100;
frog_bram[1428] = 6'b001100;
frog_bram[1429] = 6'b001100;
frog_bram[1430] = 6'b001100;
frog_bram[1431] = 6'b000000;
frog_bram[1432] = 6'b001000;
frog_bram[1433] = 6'b001100;
frog_bram[1434] = 6'b001000;
frog_bram[1435] = 6'b000000;
frog_bram[1436] = 6'b000000;
frog_bram[1437] = 6'b000000;
frog_bram[1438] = 6'b000000;
frog_bram[1439] = 6'b000000;
frog_bram[1440] = 6'b000000;
frog_bram[1441] = 6'b000000;
frog_bram[1442] = 6'b000000;
frog_bram[1443] = 6'b000000;
frog_bram[1444] = 6'b000000;
frog_bram[1445] = 6'b000000;
frog_bram[1446] = 6'b001000;
frog_bram[1447] = 6'b001000;
frog_bram[1448] = 6'b000000;
frog_bram[1449] = 6'b001100;
frog_bram[1450] = 6'b001100;
frog_bram[1451] = 6'b001100;
frog_bram[1452] = 6'b001100;
frog_bram[1453] = 6'b001100;
frog_bram[1454] = 6'b001000;
frog_bram[1455] = 6'b001000;
frog_bram[1456] = 6'b001000;
frog_bram[1457] = 6'b001000;
frog_bram[1458] = 6'b001100;
frog_bram[1459] = 6'b001100;
frog_bram[1460] = 6'b001100;
frog_bram[1461] = 6'b001100;
frog_bram[1462] = 6'b001100;
frog_bram[1463] = 6'b000000;
frog_bram[1464] = 6'b001000;
frog_bram[1465] = 6'b001000;
frog_bram[1466] = 6'b000000;
frog_bram[1467] = 6'b000000;
frog_bram[1468] = 6'b000000;
frog_bram[1469] = 6'b000000;
frog_bram[1470] = 6'b000000;
frog_bram[1471] = 6'b000000;
frog_bram[1472] = 6'b000000;
frog_bram[1473] = 6'b000000;
frog_bram[1474] = 6'b000000;
frog_bram[1475] = 6'b000000;
frog_bram[1476] = 6'b000000;
frog_bram[1477] = 6'b000000;
frog_bram[1478] = 6'b000000;
frog_bram[1479] = 6'b000000;
frog_bram[1480] = 6'b001000;
frog_bram[1481] = 6'b001100;
frog_bram[1482] = 6'b001100;
frog_bram[1483] = 6'b001100;
frog_bram[1484] = 6'b001100;
frog_bram[1485] = 6'b001000;
frog_bram[1486] = 6'b001000;
frog_bram[1487] = 6'b001000;
frog_bram[1488] = 6'b001000;
frog_bram[1489] = 6'b001000;
frog_bram[1490] = 6'b001000;
frog_bram[1491] = 6'b001100;
frog_bram[1492] = 6'b001100;
frog_bram[1493] = 6'b001100;
frog_bram[1494] = 6'b001100;
frog_bram[1495] = 6'b001000;
frog_bram[1496] = 6'b000000;
frog_bram[1497] = 6'b000000;
frog_bram[1498] = 6'b000000;
frog_bram[1499] = 6'b000000;
frog_bram[1500] = 6'b000000;
frog_bram[1501] = 6'b000000;
frog_bram[1502] = 6'b000000;
frog_bram[1503] = 6'b000000;
frog_bram[1504] = 6'b000000;
frog_bram[1505] = 6'b000000;
frog_bram[1506] = 6'b000000;
frog_bram[1507] = 6'b000000;
frog_bram[1508] = 6'b000000;
frog_bram[1509] = 6'b000000;
frog_bram[1510] = 6'b000000;
frog_bram[1511] = 6'b001000;
frog_bram[1512] = 6'b000000;
frog_bram[1513] = 6'b001100;
frog_bram[1514] = 6'b001100;
frog_bram[1515] = 6'b001100;
frog_bram[1516] = 6'b001100;
frog_bram[1517] = 6'b001100;
frog_bram[1518] = 6'b001000;
frog_bram[1519] = 6'b001000;
frog_bram[1520] = 6'b001000;
frog_bram[1521] = 6'b001000;
frog_bram[1522] = 6'b001100;
frog_bram[1523] = 6'b001100;
frog_bram[1524] = 6'b001100;
frog_bram[1525] = 6'b001100;
frog_bram[1526] = 6'b001100;
frog_bram[1527] = 6'b000000;
frog_bram[1528] = 6'b001000;
frog_bram[1529] = 6'b000000;
frog_bram[1530] = 6'b000000;
frog_bram[1531] = 6'b000000;
frog_bram[1532] = 6'b000000;
frog_bram[1533] = 6'b000000;
frog_bram[1534] = 6'b000000;
frog_bram[1535] = 6'b000000;
frog_bram[1536] = 6'b000000;
frog_bram[1537] = 6'b000000;
frog_bram[1538] = 6'b000000;
frog_bram[1539] = 6'b000000;
frog_bram[1540] = 6'b000000;
frog_bram[1541] = 6'b000000;
frog_bram[1542] = 6'b001000;
frog_bram[1543] = 6'b001100;
frog_bram[1544] = 6'b000000;
frog_bram[1545] = 6'b001100;
frog_bram[1546] = 6'b001100;
frog_bram[1547] = 6'b001100;
frog_bram[1548] = 6'b001100;
frog_bram[1549] = 6'b001100;
frog_bram[1550] = 6'b001100;
frog_bram[1551] = 6'b001000;
frog_bram[1552] = 6'b001000;
frog_bram[1553] = 6'b001100;
frog_bram[1554] = 6'b001100;
frog_bram[1555] = 6'b001100;
frog_bram[1556] = 6'b001100;
frog_bram[1557] = 6'b001100;
frog_bram[1558] = 6'b001100;
frog_bram[1559] = 6'b000000;
frog_bram[1560] = 6'b001100;
frog_bram[1561] = 6'b001000;
frog_bram[1562] = 6'b000000;
frog_bram[1563] = 6'b000000;
frog_bram[1564] = 6'b000000;
frog_bram[1565] = 6'b000000;
frog_bram[1566] = 6'b000000;
frog_bram[1567] = 6'b000000;
frog_bram[1568] = 6'b000000;
frog_bram[1569] = 6'b000000;
frog_bram[1570] = 6'b000000;
frog_bram[1571] = 6'b000000;
frog_bram[1572] = 6'b001000;
frog_bram[1573] = 6'b001000;
frog_bram[1574] = 6'b001000;
frog_bram[1575] = 6'b001000;
frog_bram[1576] = 6'b001100;
frog_bram[1577] = 6'b001000;
frog_bram[1578] = 6'b001100;
frog_bram[1579] = 6'b001100;
frog_bram[1580] = 6'b001100;
frog_bram[1581] = 6'b001100;
frog_bram[1582] = 6'b001100;
frog_bram[1583] = 6'b001000;
frog_bram[1584] = 6'b001000;
frog_bram[1585] = 6'b001100;
frog_bram[1586] = 6'b001100;
frog_bram[1587] = 6'b001100;
frog_bram[1588] = 6'b001100;
frog_bram[1589] = 6'b001100;
frog_bram[1590] = 6'b001000;
frog_bram[1591] = 6'b001100;
frog_bram[1592] = 6'b001000;
frog_bram[1593] = 6'b001000;
frog_bram[1594] = 6'b001000;
frog_bram[1595] = 6'b001000;
frog_bram[1596] = 6'b000000;
frog_bram[1597] = 6'b000000;
frog_bram[1598] = 6'b000000;
frog_bram[1599] = 6'b000000;
frog_bram[1600] = 6'b000000;
frog_bram[1601] = 6'b000000;
frog_bram[1602] = 6'b000000;
frog_bram[1603] = 6'b001000;
frog_bram[1604] = 6'b001000;
frog_bram[1605] = 6'b001000;
frog_bram[1606] = 6'b001000;
frog_bram[1607] = 6'b001000;
frog_bram[1608] = 6'b001000;
frog_bram[1609] = 6'b000000;
frog_bram[1610] = 6'b001000;
frog_bram[1611] = 6'b001100;
frog_bram[1612] = 6'b001100;
frog_bram[1613] = 6'b001100;
frog_bram[1614] = 6'b001000;
frog_bram[1615] = 6'b001000;
frog_bram[1616] = 6'b001000;
frog_bram[1617] = 6'b001000;
frog_bram[1618] = 6'b001100;
frog_bram[1619] = 6'b001100;
frog_bram[1620] = 6'b001100;
frog_bram[1621] = 6'b001000;
frog_bram[1622] = 6'b000000;
frog_bram[1623] = 6'b001000;
frog_bram[1624] = 6'b001000;
frog_bram[1625] = 6'b001000;
frog_bram[1626] = 6'b001000;
frog_bram[1627] = 6'b001000;
frog_bram[1628] = 6'b001000;
frog_bram[1629] = 6'b000000;
frog_bram[1630] = 6'b000000;
frog_bram[1631] = 6'b000000;
frog_bram[1632] = 6'b000000;
frog_bram[1633] = 6'b000000;
frog_bram[1634] = 6'b001100;
frog_bram[1635] = 6'b001100;
frog_bram[1636] = 6'b001100;
frog_bram[1637] = 6'b001000;
frog_bram[1638] = 6'b001000;
frog_bram[1639] = 6'b001000;
frog_bram[1640] = 6'b000000;
frog_bram[1641] = 6'b000000;
frog_bram[1642] = 6'b001000;
frog_bram[1643] = 6'b001100;
frog_bram[1644] = 6'b001100;
frog_bram[1645] = 6'b001100;
frog_bram[1646] = 6'b001100;
frog_bram[1647] = 6'b001100;
frog_bram[1648] = 6'b001100;
frog_bram[1649] = 6'b001100;
frog_bram[1650] = 6'b001100;
frog_bram[1651] = 6'b001100;
frog_bram[1652] = 6'b001100;
frog_bram[1653] = 6'b001000;
frog_bram[1654] = 6'b000000;
frog_bram[1655] = 6'b000000;
frog_bram[1656] = 6'b001000;
frog_bram[1657] = 6'b001000;
frog_bram[1658] = 6'b001000;
frog_bram[1659] = 6'b001100;
frog_bram[1660] = 6'b001100;
frog_bram[1661] = 6'b001100;
frog_bram[1662] = 6'b000000;
frog_bram[1663] = 6'b000000;
frog_bram[1664] = 6'b000000;
frog_bram[1665] = 6'b000000;
frog_bram[1666] = 6'b001100;
frog_bram[1667] = 6'b001100;
frog_bram[1668] = 6'b001100;
frog_bram[1669] = 6'b001000;
frog_bram[1670] = 6'b000000;
frog_bram[1671] = 6'b000000;
frog_bram[1672] = 6'b000000;
frog_bram[1673] = 6'b001100;
frog_bram[1674] = 6'b001100;
frog_bram[1675] = 6'b001100;
frog_bram[1676] = 6'b001100;
frog_bram[1677] = 6'b001100;
frog_bram[1678] = 6'b001100;
frog_bram[1679] = 6'b001100;
frog_bram[1680] = 6'b001100;
frog_bram[1681] = 6'b001100;
frog_bram[1682] = 6'b001100;
frog_bram[1683] = 6'b001100;
frog_bram[1684] = 6'b001100;
frog_bram[1685] = 6'b001100;
frog_bram[1686] = 6'b001100;
frog_bram[1687] = 6'b000000;
frog_bram[1688] = 6'b000000;
frog_bram[1689] = 6'b000000;
frog_bram[1690] = 6'b001000;
frog_bram[1691] = 6'b001100;
frog_bram[1692] = 6'b001100;
frog_bram[1693] = 6'b001100;
frog_bram[1694] = 6'b000000;
frog_bram[1695] = 6'b000000;
frog_bram[1696] = 6'b000000;
frog_bram[1697] = 6'b000000;
frog_bram[1698] = 6'b001100;
frog_bram[1699] = 6'b001100;
frog_bram[1700] = 6'b001100;
frog_bram[1701] = 6'b000000;
frog_bram[1702] = 6'b000000;
frog_bram[1703] = 6'b000000;
frog_bram[1704] = 6'b001100;
frog_bram[1705] = 6'b001100;
frog_bram[1706] = 6'b001100;
frog_bram[1707] = 6'b001000;
frog_bram[1708] = 6'b001000;
frog_bram[1709] = 6'b001000;
frog_bram[1710] = 6'b001100;
frog_bram[1711] = 6'b001100;
frog_bram[1712] = 6'b001100;
frog_bram[1713] = 6'b001100;
frog_bram[1714] = 6'b001100;
frog_bram[1715] = 6'b001100;
frog_bram[1716] = 6'b001100;
frog_bram[1717] = 6'b001100;
frog_bram[1718] = 6'b001100;
frog_bram[1719] = 6'b001100;
frog_bram[1720] = 6'b000000;
frog_bram[1721] = 6'b000000;
frog_bram[1722] = 6'b000000;
frog_bram[1723] = 6'b001100;
frog_bram[1724] = 6'b001100;
frog_bram[1725] = 6'b001100;
frog_bram[1726] = 6'b000000;
frog_bram[1727] = 6'b000000;
frog_bram[1728] = 6'b000000;
frog_bram[1729] = 6'b000000;
frog_bram[1730] = 6'b001100;
frog_bram[1731] = 6'b001100;
frog_bram[1732] = 6'b001100;
frog_bram[1733] = 6'b001100;
frog_bram[1734] = 6'b000000;
frog_bram[1735] = 6'b000000;
frog_bram[1736] = 6'b001100;
frog_bram[1737] = 6'b001100;
frog_bram[1738] = 6'b001000;
frog_bram[1739] = 6'b110000;
frog_bram[1740] = 6'b110000;
frog_bram[1741] = 6'b001000;
frog_bram[1742] = 6'b001000;
frog_bram[1743] = 6'b001100;
frog_bram[1744] = 6'b001100;
frog_bram[1745] = 6'b001100;
frog_bram[1746] = 6'b001100;
frog_bram[1747] = 6'b110000;
frog_bram[1748] = 6'b110000;
frog_bram[1749] = 6'b001100;
frog_bram[1750] = 6'b001100;
frog_bram[1751] = 6'b001100;
frog_bram[1752] = 6'b000000;
frog_bram[1753] = 6'b000000;
frog_bram[1754] = 6'b001100;
frog_bram[1755] = 6'b001100;
frog_bram[1756] = 6'b001100;
frog_bram[1757] = 6'b001100;
frog_bram[1758] = 6'b000000;
frog_bram[1759] = 6'b000000;
frog_bram[1760] = 6'b000000;
frog_bram[1761] = 6'b000000;
frog_bram[1762] = 6'b001100;
frog_bram[1763] = 6'b001100;
frog_bram[1764] = 6'b001100;
frog_bram[1765] = 6'b001100;
frog_bram[1766] = 6'b001000;
frog_bram[1767] = 6'b000000;
frog_bram[1768] = 6'b001000;
frog_bram[1769] = 6'b001000;
frog_bram[1770] = 6'b100000;
frog_bram[1771] = 6'b010000;
frog_bram[1772] = 6'b010000;
frog_bram[1773] = 6'b110000;
frog_bram[1774] = 6'b001000;
frog_bram[1775] = 6'b001100;
frog_bram[1776] = 6'b001100;
frog_bram[1777] = 6'b001100;
frog_bram[1778] = 6'b110000;
frog_bram[1779] = 6'b010000;
frog_bram[1780] = 6'b010000;
frog_bram[1781] = 6'b110000;
frog_bram[1782] = 6'b001100;
frog_bram[1783] = 6'b001100;
frog_bram[1784] = 6'b000000;
frog_bram[1785] = 6'b001000;
frog_bram[1786] = 6'b001100;
frog_bram[1787] = 6'b001100;
frog_bram[1788] = 6'b001100;
frog_bram[1789] = 6'b001100;
frog_bram[1790] = 6'b000000;
frog_bram[1791] = 6'b000000;
frog_bram[1792] = 6'b000000;
frog_bram[1793] = 6'b000000;
frog_bram[1794] = 6'b001100;
frog_bram[1795] = 6'b001100;
frog_bram[1796] = 6'b001100;
frog_bram[1797] = 6'b000100;
frog_bram[1798] = 6'b001000;
frog_bram[1799] = 6'b000000;
frog_bram[1800] = 6'b000000;
frog_bram[1801] = 6'b001000;
frog_bram[1802] = 6'b110000;
frog_bram[1803] = 6'b010000;
frog_bram[1804] = 6'b010000;
frog_bram[1805] = 6'b110000;
frog_bram[1806] = 6'b001000;
frog_bram[1807] = 6'b001100;
frog_bram[1808] = 6'b001100;
frog_bram[1809] = 6'b001100;
frog_bram[1810] = 6'b110000;
frog_bram[1811] = 6'b010000;
frog_bram[1812] = 6'b010000;
frog_bram[1813] = 6'b110000;
frog_bram[1814] = 6'b001100;
frog_bram[1815] = 6'b001100;
frog_bram[1816] = 6'b000000;
frog_bram[1817] = 6'b000100;
frog_bram[1818] = 6'b000100;
frog_bram[1819] = 6'b001100;
frog_bram[1820] = 6'b001100;
frog_bram[1821] = 6'b001100;
frog_bram[1822] = 6'b000000;
frog_bram[1823] = 6'b000000;
frog_bram[1824] = 6'b000000;
frog_bram[1825] = 6'b000000;
frog_bram[1826] = 6'b000000;
frog_bram[1827] = 6'b001100;
frog_bram[1828] = 6'b001000;
frog_bram[1829] = 6'b001000;
frog_bram[1830] = 6'b000000;
frog_bram[1831] = 6'b000000;
frog_bram[1832] = 6'b000000;
frog_bram[1833] = 6'b001000;
frog_bram[1834] = 6'b001000;
frog_bram[1835] = 6'b110000;
frog_bram[1836] = 6'b110000;
frog_bram[1837] = 6'b001000;
frog_bram[1838] = 6'b001100;
frog_bram[1839] = 6'b001100;
frog_bram[1840] = 6'b001100;
frog_bram[1841] = 6'b001100;
frog_bram[1842] = 6'b001100;
frog_bram[1843] = 6'b110000;
frog_bram[1844] = 6'b110000;
frog_bram[1845] = 6'b001100;
frog_bram[1846] = 6'b001100;
frog_bram[1847] = 6'b000000;
frog_bram[1848] = 6'b000000;
frog_bram[1849] = 6'b000000;
frog_bram[1850] = 6'b001000;
frog_bram[1851] = 6'b001000;
frog_bram[1852] = 6'b001100;
frog_bram[1853] = 6'b000000;
frog_bram[1854] = 6'b000000;
frog_bram[1855] = 6'b000000;
frog_bram[1856] = 6'b000000;
frog_bram[1857] = 6'b000000;
frog_bram[1858] = 6'b000000;
frog_bram[1859] = 6'b001100;
frog_bram[1860] = 6'b000100;
frog_bram[1861] = 6'b001100;
frog_bram[1862] = 6'b001100;
frog_bram[1863] = 6'b000000;
frog_bram[1864] = 6'b000000;
frog_bram[1865] = 6'b000000;
frog_bram[1866] = 6'b001000;
frog_bram[1867] = 6'b001000;
frog_bram[1868] = 6'b001000;
frog_bram[1869] = 6'b001100;
frog_bram[1870] = 6'b001100;
frog_bram[1871] = 6'b001100;
frog_bram[1872] = 6'b001100;
frog_bram[1873] = 6'b001100;
frog_bram[1874] = 6'b001100;
frog_bram[1875] = 6'b001100;
frog_bram[1876] = 6'b001100;
frog_bram[1877] = 6'b001000;
frog_bram[1878] = 6'b000000;
frog_bram[1879] = 6'b000000;
frog_bram[1880] = 6'b000000;
frog_bram[1881] = 6'b001100;
frog_bram[1882] = 6'b001100;
frog_bram[1883] = 6'b000100;
frog_bram[1884] = 6'b001100;
frog_bram[1885] = 6'b000000;
frog_bram[1886] = 6'b000000;
frog_bram[1887] = 6'b000000;
frog_bram[1888] = 6'b000000;
frog_bram[1889] = 6'b000000;
frog_bram[1890] = 6'b000000;
frog_bram[1891] = 6'b001100;
frog_bram[1892] = 6'b001000;
frog_bram[1893] = 6'b000000;
frog_bram[1894] = 6'b001100;
frog_bram[1895] = 6'b001000;
frog_bram[1896] = 6'b000000;
frog_bram[1897] = 6'b000000;
frog_bram[1898] = 6'b000000;
frog_bram[1899] = 6'b001000;
frog_bram[1900] = 6'b001100;
frog_bram[1901] = 6'b001100;
frog_bram[1902] = 6'b001100;
frog_bram[1903] = 6'b001100;
frog_bram[1904] = 6'b001100;
frog_bram[1905] = 6'b001100;
frog_bram[1906] = 6'b001100;
frog_bram[1907] = 6'b001100;
frog_bram[1908] = 6'b001000;
frog_bram[1909] = 6'b000000;
frog_bram[1910] = 6'b000000;
frog_bram[1911] = 6'b000000;
frog_bram[1912] = 6'b001000;
frog_bram[1913] = 6'b001100;
frog_bram[1914] = 6'b000000;
frog_bram[1915] = 6'b001000;
frog_bram[1916] = 6'b001100;
frog_bram[1917] = 6'b000000;
frog_bram[1918] = 6'b000000;
frog_bram[1919] = 6'b000000;
frog_bram[1920] = 6'b000000;
frog_bram[1921] = 6'b000000;
frog_bram[1922] = 6'b000000;
frog_bram[1923] = 6'b001100;
frog_bram[1924] = 6'b001000;
frog_bram[1925] = 6'b000000;
frog_bram[1926] = 6'b001000;
frog_bram[1927] = 6'b001000;
frog_bram[1928] = 6'b000000;
frog_bram[1929] = 6'b000000;
frog_bram[1930] = 6'b000000;
frog_bram[1931] = 6'b000000;
frog_bram[1932] = 6'b001100;
frog_bram[1933] = 6'b001100;
frog_bram[1934] = 6'b000100;
frog_bram[1935] = 6'b001100;
frog_bram[1936] = 6'b001100;
frog_bram[1937] = 6'b000100;
frog_bram[1938] = 6'b001100;
frog_bram[1939] = 6'b001100;
frog_bram[1940] = 6'b000000;
frog_bram[1941] = 6'b000000;
frog_bram[1942] = 6'b000000;
frog_bram[1943] = 6'b000000;
frog_bram[1944] = 6'b001000;
frog_bram[1945] = 6'b001000;
frog_bram[1946] = 6'b000000;
frog_bram[1947] = 6'b001000;
frog_bram[1948] = 6'b001100;
frog_bram[1949] = 6'b000000;
frog_bram[1950] = 6'b000000;
frog_bram[1951] = 6'b000000;
frog_bram[1952] = 6'b000000;
frog_bram[1953] = 6'b000000;
frog_bram[1954] = 6'b000000;
frog_bram[1955] = 6'b000000;
frog_bram[1956] = 6'b000000;
frog_bram[1957] = 6'b000000;
frog_bram[1958] = 6'b000000;
frog_bram[1959] = 6'b000000;
frog_bram[1960] = 6'b000000;
frog_bram[1961] = 6'b000000;
frog_bram[1962] = 6'b000000;
frog_bram[1963] = 6'b000000;
frog_bram[1964] = 6'b000000;
frog_bram[1965] = 6'b001000;
frog_bram[1966] = 6'b001000;
frog_bram[1967] = 6'b001100;
frog_bram[1968] = 6'b001100;
frog_bram[1969] = 6'b001000;
frog_bram[1970] = 6'b001000;
frog_bram[1971] = 6'b000000;
frog_bram[1972] = 6'b000000;
frog_bram[1973] = 6'b000000;
frog_bram[1974] = 6'b000000;
frog_bram[1975] = 6'b000000;
frog_bram[1976] = 6'b000000;
frog_bram[1977] = 6'b000000;
frog_bram[1978] = 6'b000000;
frog_bram[1979] = 6'b000000;
frog_bram[1980] = 6'b000000;
frog_bram[1981] = 6'b000000;
frog_bram[1982] = 6'b000000;
frog_bram[1983] = 6'b000000;
frog_bram[1984] = 6'b000000;
frog_bram[1985] = 6'b000000;
frog_bram[1986] = 6'b000000;
frog_bram[1987] = 6'b000000;
frog_bram[1988] = 6'b000000;
frog_bram[1989] = 6'b000000;
frog_bram[1990] = 6'b000000;
frog_bram[1991] = 6'b000000;
frog_bram[1992] = 6'b000000;
frog_bram[1993] = 6'b000000;
frog_bram[1994] = 6'b000000;
frog_bram[1995] = 6'b000000;
frog_bram[1996] = 6'b000000;
frog_bram[1997] = 6'b000000;
frog_bram[1998] = 6'b000000;
frog_bram[1999] = 6'b000000;
frog_bram[2000] = 6'b000000;
frog_bram[2001] = 6'b000000;
frog_bram[2002] = 6'b000000;
frog_bram[2003] = 6'b000000;
frog_bram[2004] = 6'b000000;
frog_bram[2005] = 6'b000000;
frog_bram[2006] = 6'b000000;
frog_bram[2007] = 6'b000000;
frog_bram[2008] = 6'b000000;
frog_bram[2009] = 6'b000000;
frog_bram[2010] = 6'b000000;
frog_bram[2011] = 6'b000000;
frog_bram[2012] = 6'b000000;
frog_bram[2013] = 6'b000000;
frog_bram[2014] = 6'b000000;
frog_bram[2015] = 6'b000000;
frog_bram[2016] = 6'b000000;
frog_bram[2017] = 6'b000000;
frog_bram[2018] = 6'b000000;
frog_bram[2019] = 6'b000000;
frog_bram[2020] = 6'b000000;
frog_bram[2021] = 6'b000000;
frog_bram[2022] = 6'b000000;
frog_bram[2023] = 6'b000000;
frog_bram[2024] = 6'b000000;
frog_bram[2025] = 6'b000000;
frog_bram[2026] = 6'b000000;
frog_bram[2027] = 6'b000000;
frog_bram[2028] = 6'b000000;
frog_bram[2029] = 6'b000000;
frog_bram[2030] = 6'b000000;
frog_bram[2031] = 6'b000000;
frog_bram[2032] = 6'b000000;
frog_bram[2033] = 6'b000000;
frog_bram[2034] = 6'b000000;
frog_bram[2035] = 6'b000000;
frog_bram[2036] = 6'b000000;
frog_bram[2037] = 6'b000000;
frog_bram[2038] = 6'b000000;
frog_bram[2039] = 6'b000000;
frog_bram[2040] = 6'b000000;
frog_bram[2041] = 6'b000000;
frog_bram[2042] = 6'b000000;
frog_bram[2043] = 6'b000000;
frog_bram[2044] = 6'b000000;
frog_bram[2045] = 6'b000000;
frog_bram[2046] = 6'b000000;
frog_bram[2047] = 6'b000000;
        // Add more initialization here for the left-facing sprite (2048 - 3071)
frog_bram[2048] = 6'b000000;
frog_bram[2049] = 6'b000000;
frog_bram[2050] = 6'b000000;
frog_bram[2051] = 6'b000000;
frog_bram[2052] = 6'b000000;
frog_bram[2053] = 6'b000000;
frog_bram[2054] = 6'b000000;
frog_bram[2055] = 6'b000000;
frog_bram[2056] = 6'b000000;
frog_bram[2057] = 6'b000000;
frog_bram[2058] = 6'b000000;
frog_bram[2059] = 6'b000000;
frog_bram[2060] = 6'b000000;
frog_bram[2061] = 6'b000000;
frog_bram[2062] = 6'b000000;
frog_bram[2063] = 6'b000000;
frog_bram[2064] = 6'b000000;
frog_bram[2065] = 6'b000000;
frog_bram[2066] = 6'b000000;
frog_bram[2067] = 6'b000000;
frog_bram[2068] = 6'b000000;
frog_bram[2069] = 6'b000000;
frog_bram[2070] = 6'b000000;
frog_bram[2071] = 6'b000000;
frog_bram[2072] = 6'b001000;
frog_bram[2073] = 6'b001100;
frog_bram[2074] = 6'b000000;
frog_bram[2075] = 6'b001000;
frog_bram[2076] = 6'b001100;
frog_bram[2077] = 6'b000000;
frog_bram[2078] = 6'b000000;
frog_bram[2079] = 6'b000000;
frog_bram[2080] = 6'b000000;
frog_bram[2081] = 6'b000000;
frog_bram[2082] = 6'b000000;
frog_bram[2083] = 6'b000000;
frog_bram[2084] = 6'b000000;
frog_bram[2085] = 6'b000000;
frog_bram[2086] = 6'b000000;
frog_bram[2087] = 6'b000000;
frog_bram[2088] = 6'b000000;
frog_bram[2089] = 6'b000000;
frog_bram[2090] = 6'b000000;
frog_bram[2091] = 6'b000000;
frog_bram[2092] = 6'b000000;
frog_bram[2093] = 6'b000000;
frog_bram[2094] = 6'b000000;
frog_bram[2095] = 6'b000000;
frog_bram[2096] = 6'b000000;
frog_bram[2097] = 6'b000000;
frog_bram[2098] = 6'b000000;
frog_bram[2099] = 6'b000000;
frog_bram[2100] = 6'b000000;
frog_bram[2101] = 6'b000000;
frog_bram[2102] = 6'b000000;
frog_bram[2103] = 6'b000000;
frog_bram[2104] = 6'b001000;
frog_bram[2105] = 6'b001100;
frog_bram[2106] = 6'b001100;
frog_bram[2107] = 6'b001100;
frog_bram[2108] = 6'b001100;
frog_bram[2109] = 6'b000000;
frog_bram[2110] = 6'b000000;
frog_bram[2111] = 6'b000000;
frog_bram[2112] = 6'b000000;
frog_bram[2113] = 6'b000000;
frog_bram[2114] = 6'b000000;
frog_bram[2115] = 6'b000000;
frog_bram[2116] = 6'b000000;
frog_bram[2117] = 6'b000000;
frog_bram[2118] = 6'b000000;
frog_bram[2119] = 6'b001100;
frog_bram[2120] = 6'b001100;
frog_bram[2121] = 6'b001100;
frog_bram[2122] = 6'b001100;
frog_bram[2123] = 6'b001100;
frog_bram[2124] = 6'b001100;
frog_bram[2125] = 6'b000000;
frog_bram[2126] = 6'b000000;
frog_bram[2127] = 6'b000000;
frog_bram[2128] = 6'b000000;
frog_bram[2129] = 6'b000000;
frog_bram[2130] = 6'b000000;
frog_bram[2131] = 6'b000000;
frog_bram[2132] = 6'b000000;
frog_bram[2133] = 6'b000000;
frog_bram[2134] = 6'b001000;
frog_bram[2135] = 6'b001100;
frog_bram[2136] = 6'b000100;
frog_bram[2137] = 6'b001000;
frog_bram[2138] = 6'b001100;
frog_bram[2139] = 6'b001100;
frog_bram[2140] = 6'b001100;
frog_bram[2141] = 6'b001000;
frog_bram[2142] = 6'b000000;
frog_bram[2143] = 6'b000000;
frog_bram[2144] = 6'b000000;
frog_bram[2145] = 6'b000000;
frog_bram[2146] = 6'b000000;
frog_bram[2147] = 6'b001100;
frog_bram[2148] = 6'b001100;
frog_bram[2149] = 6'b001100;
frog_bram[2150] = 6'b001100;
frog_bram[2151] = 6'b001100;
frog_bram[2152] = 6'b001100;
frog_bram[2153] = 6'b001100;
frog_bram[2154] = 6'b001100;
frog_bram[2155] = 6'b001100;
frog_bram[2156] = 6'b001100;
frog_bram[2157] = 6'b001000;
frog_bram[2158] = 6'b000000;
frog_bram[2159] = 6'b000000;
frog_bram[2160] = 6'b000000;
frog_bram[2161] = 6'b000000;
frog_bram[2162] = 6'b000000;
frog_bram[2163] = 6'b000000;
frog_bram[2164] = 6'b000000;
frog_bram[2165] = 6'b000000;
frog_bram[2166] = 6'b001000;
frog_bram[2167] = 6'b001100;
frog_bram[2168] = 6'b001100;
frog_bram[2169] = 6'b001100;
frog_bram[2170] = 6'b001100;
frog_bram[2171] = 6'b001100;
frog_bram[2172] = 6'b001100;
frog_bram[2173] = 6'b001000;
frog_bram[2174] = 6'b000000;
frog_bram[2175] = 6'b000000;
frog_bram[2176] = 6'b000000;
frog_bram[2177] = 6'b000000;
frog_bram[2178] = 6'b000000;
frog_bram[2179] = 6'b001000;
frog_bram[2180] = 6'b001000;
frog_bram[2181] = 6'b000100;
frog_bram[2182] = 6'b001000;
frog_bram[2183] = 6'b001100;
frog_bram[2184] = 6'b001100;
frog_bram[2185] = 6'b001100;
frog_bram[2186] = 6'b001100;
frog_bram[2187] = 6'b001100;
frog_bram[2188] = 6'b001100;
frog_bram[2189] = 6'b001000;
frog_bram[2190] = 6'b001000;
frog_bram[2191] = 6'b000000;
frog_bram[2192] = 6'b000000;
frog_bram[2193] = 6'b000000;
frog_bram[2194] = 6'b000000;
frog_bram[2195] = 6'b000000;
frog_bram[2196] = 6'b000000;
frog_bram[2197] = 6'b000000;
frog_bram[2198] = 6'b000000;
frog_bram[2199] = 6'b000000;
frog_bram[2200] = 6'b000000;
frog_bram[2201] = 6'b001000;
frog_bram[2202] = 6'b001100;
frog_bram[2203] = 6'b001100;
frog_bram[2204] = 6'b001100;
frog_bram[2205] = 6'b001000;
frog_bram[2206] = 6'b000000;
frog_bram[2207] = 6'b000000;
frog_bram[2208] = 6'b000000;
frog_bram[2209] = 6'b000000;
frog_bram[2210] = 6'b000000;
frog_bram[2211] = 6'b000000;
frog_bram[2212] = 6'b000000;
frog_bram[2213] = 6'b001100;
frog_bram[2214] = 6'b001000;
frog_bram[2215] = 6'b000100;
frog_bram[2216] = 6'b001100;
frog_bram[2217] = 6'b001100;
frog_bram[2218] = 6'b000000;
frog_bram[2219] = 6'b001000;
frog_bram[2220] = 6'b001000;
frog_bram[2221] = 6'b001000;
frog_bram[2222] = 6'b001000;
frog_bram[2223] = 6'b000000;
frog_bram[2224] = 6'b000000;
frog_bram[2225] = 6'b000000;
frog_bram[2226] = 6'b000000;
frog_bram[2227] = 6'b001000;
frog_bram[2228] = 6'b001000;
frog_bram[2229] = 6'b001000;
frog_bram[2230] = 6'b001000;
frog_bram[2231] = 6'b001000;
frog_bram[2232] = 6'b001000;
frog_bram[2233] = 6'b000000;
frog_bram[2234] = 6'b001000;
frog_bram[2235] = 6'b001100;
frog_bram[2236] = 6'b001100;
frog_bram[2237] = 6'b001100;
frog_bram[2238] = 6'b001000;
frog_bram[2239] = 6'b000000;
frog_bram[2240] = 6'b000000;
frog_bram[2241] = 6'b000000;
frog_bram[2242] = 6'b000000;
frog_bram[2243] = 6'b001000;
frog_bram[2244] = 6'b001100;
frog_bram[2245] = 6'b001100;
frog_bram[2246] = 6'b000000;
frog_bram[2247] = 6'b000100;
frog_bram[2248] = 6'b001000;
frog_bram[2249] = 6'b000000;
frog_bram[2250] = 6'b000000;
frog_bram[2251] = 6'b000000;
frog_bram[2252] = 6'b001000;
frog_bram[2253] = 6'b001000;
frog_bram[2254] = 6'b001000;
frog_bram[2255] = 6'b001000;
frog_bram[2256] = 6'b000000;
frog_bram[2257] = 6'b000000;
frog_bram[2258] = 6'b001000;
frog_bram[2259] = 6'b001100;
frog_bram[2260] = 6'b001100;
frog_bram[2261] = 6'b001100;
frog_bram[2262] = 6'b001100;
frog_bram[2263] = 6'b001100;
frog_bram[2264] = 6'b001000;
frog_bram[2265] = 6'b001000;
frog_bram[2266] = 6'b000000;
frog_bram[2267] = 6'b001100;
frog_bram[2268] = 6'b001100;
frog_bram[2269] = 6'b001100;
frog_bram[2270] = 6'b001000;
frog_bram[2271] = 6'b000000;
frog_bram[2272] = 6'b000000;
frog_bram[2273] = 6'b000000;
frog_bram[2274] = 6'b000000;
frog_bram[2275] = 6'b001000;
frog_bram[2276] = 6'b001000;
frog_bram[2277] = 6'b000000;
frog_bram[2278] = 6'b000000;
frog_bram[2279] = 6'b000000;
frog_bram[2280] = 6'b000000;
frog_bram[2281] = 6'b000000;
frog_bram[2282] = 6'b000000;
frog_bram[2283] = 6'b000000;
frog_bram[2284] = 6'b001000;
frog_bram[2285] = 6'b001000;
frog_bram[2286] = 6'b001000;
frog_bram[2287] = 6'b001100;
frog_bram[2288] = 6'b001000;
frog_bram[2289] = 6'b000000;
frog_bram[2290] = 6'b001000;
frog_bram[2291] = 6'b001000;
frog_bram[2292] = 6'b001000;
frog_bram[2293] = 6'b001000;
frog_bram[2294] = 6'b001100;
frog_bram[2295] = 6'b001100;
frog_bram[2296] = 6'b001100;
frog_bram[2297] = 6'b001100;
frog_bram[2298] = 6'b001100;
frog_bram[2299] = 6'b001100;
frog_bram[2300] = 6'b001100;
frog_bram[2301] = 6'b001100;
frog_bram[2302] = 6'b000000;
frog_bram[2303] = 6'b000000;
frog_bram[2304] = 6'b000000;
frog_bram[2305] = 6'b000000;
frog_bram[2306] = 6'b000000;
frog_bram[2307] = 6'b000000;
frog_bram[2308] = 6'b000000;
frog_bram[2309] = 6'b000000;
frog_bram[2310] = 6'b000000;
frog_bram[2311] = 6'b001100;
frog_bram[2312] = 6'b001100;
frog_bram[2313] = 6'b001100;
frog_bram[2314] = 6'b001100;
frog_bram[2315] = 6'b000000;
frog_bram[2316] = 6'b000000;
frog_bram[2317] = 6'b001000;
frog_bram[2318] = 6'b001100;
frog_bram[2319] = 6'b000000;
frog_bram[2320] = 6'b000000;
frog_bram[2321] = 6'b001000;
frog_bram[2322] = 6'b000000;
frog_bram[2323] = 6'b000000;
frog_bram[2324] = 6'b000000;
frog_bram[2325] = 6'b000000;
frog_bram[2326] = 6'b001000;
frog_bram[2327] = 6'b001000;
frog_bram[2328] = 6'b001000;
frog_bram[2329] = 6'b001100;
frog_bram[2330] = 6'b001100;
frog_bram[2331] = 6'b001100;
frog_bram[2332] = 6'b001100;
frog_bram[2333] = 6'b001000;
frog_bram[2334] = 6'b000000;
frog_bram[2335] = 6'b000000;
frog_bram[2336] = 6'b000000;
frog_bram[2337] = 6'b000000;
frog_bram[2338] = 6'b000000;
frog_bram[2339] = 6'b000000;
frog_bram[2340] = 6'b000000;
frog_bram[2341] = 6'b000000;
frog_bram[2342] = 6'b001100;
frog_bram[2343] = 6'b001100;
frog_bram[2344] = 6'b001100;
frog_bram[2345] = 6'b001100;
frog_bram[2346] = 6'b001100;
frog_bram[2347] = 6'b001100;
frog_bram[2348] = 6'b000000;
frog_bram[2349] = 6'b000000;
frog_bram[2350] = 6'b001000;
frog_bram[2351] = 6'b001100;
frog_bram[2352] = 6'b001100;
frog_bram[2353] = 6'b001100;
frog_bram[2354] = 6'b001100;
frog_bram[2355] = 6'b001100;
frog_bram[2356] = 6'b001000;
frog_bram[2357] = 6'b001000;
frog_bram[2358] = 6'b000000;
frog_bram[2359] = 6'b000000;
frog_bram[2360] = 6'b000000;
frog_bram[2361] = 6'b001000;
frog_bram[2362] = 6'b001000;
frog_bram[2363] = 6'b001000;
frog_bram[2364] = 6'b000000;
frog_bram[2365] = 6'b000000;
frog_bram[2366] = 6'b000000;
frog_bram[2367] = 6'b000000;
frog_bram[2368] = 6'b000000;
frog_bram[2369] = 6'b000000;
frog_bram[2370] = 6'b000000;
frog_bram[2371] = 6'b000000;
frog_bram[2372] = 6'b000000;
frog_bram[2373] = 6'b001000;
frog_bram[2374] = 6'b001100;
frog_bram[2375] = 6'b110000;
frog_bram[2376] = 6'b110000;
frog_bram[2377] = 6'b001100;
frog_bram[2378] = 6'b001100;
frog_bram[2379] = 6'b001100;
frog_bram[2380] = 6'b001000;
frog_bram[2381] = 6'b001000;
frog_bram[2382] = 6'b001100;
frog_bram[2383] = 6'b001100;
frog_bram[2384] = 6'b001100;
frog_bram[2385] = 6'b001100;
frog_bram[2386] = 6'b001100;
frog_bram[2387] = 6'b001100;
frog_bram[2388] = 6'b001100;
frog_bram[2389] = 6'b001100;
frog_bram[2390] = 6'b001000;
frog_bram[2391] = 6'b001000;
frog_bram[2392] = 6'b001000;
frog_bram[2393] = 6'b000000;
frog_bram[2394] = 6'b000000;
frog_bram[2395] = 6'b000000;
frog_bram[2396] = 6'b000000;
frog_bram[2397] = 6'b000000;
frog_bram[2398] = 6'b000000;
frog_bram[2399] = 6'b000000;
frog_bram[2400] = 6'b000000;
frog_bram[2401] = 6'b000000;
frog_bram[2402] = 6'b000000;
frog_bram[2403] = 6'b000000;
frog_bram[2404] = 6'b001000;
frog_bram[2405] = 6'b001100;
frog_bram[2406] = 6'b110000;
frog_bram[2407] = 6'b010000;
frog_bram[2408] = 6'b010000;
frog_bram[2409] = 6'b110000;
frog_bram[2410] = 6'b001100;
frog_bram[2411] = 6'b001100;
frog_bram[2412] = 6'b001100;
frog_bram[2413] = 6'b001100;
frog_bram[2414] = 6'b001100;
frog_bram[2415] = 6'b001100;
frog_bram[2416] = 6'b001100;
frog_bram[2417] = 6'b001100;
frog_bram[2418] = 6'b001100;
frog_bram[2419] = 6'b001100;
frog_bram[2420] = 6'b001100;
frog_bram[2421] = 6'b001100;
frog_bram[2422] = 6'b001000;
frog_bram[2423] = 6'b001100;
frog_bram[2424] = 6'b001100;
frog_bram[2425] = 6'b001000;
frog_bram[2426] = 6'b001000;
frog_bram[2427] = 6'b000000;
frog_bram[2428] = 6'b000000;
frog_bram[2429] = 6'b000000;
frog_bram[2430] = 6'b000000;
frog_bram[2431] = 6'b000000;
frog_bram[2432] = 6'b000000;
frog_bram[2433] = 6'b000000;
frog_bram[2434] = 6'b000000;
frog_bram[2435] = 6'b001100;
frog_bram[2436] = 6'b001100;
frog_bram[2437] = 6'b001100;
frog_bram[2438] = 6'b110000;
frog_bram[2439] = 6'b010000;
frog_bram[2440] = 6'b010000;
frog_bram[2441] = 6'b110000;
frog_bram[2442] = 6'b001100;
frog_bram[2443] = 6'b001100;
frog_bram[2444] = 6'b001100;
frog_bram[2445] = 6'b001100;
frog_bram[2446] = 6'b001100;
frog_bram[2447] = 6'b001100;
frog_bram[2448] = 6'b001100;
frog_bram[2449] = 6'b001100;
frog_bram[2450] = 6'b001100;
frog_bram[2451] = 6'b001100;
frog_bram[2452] = 6'b001100;
frog_bram[2453] = 6'b001000;
frog_bram[2454] = 6'b001000;
frog_bram[2455] = 6'b001100;
frog_bram[2456] = 6'b001100;
frog_bram[2457] = 6'b001100;
frog_bram[2458] = 6'b001000;
frog_bram[2459] = 6'b000000;
frog_bram[2460] = 6'b000000;
frog_bram[2461] = 6'b000000;
frog_bram[2462] = 6'b000000;
frog_bram[2463] = 6'b000000;
frog_bram[2464] = 6'b000000;
frog_bram[2465] = 6'b000000;
frog_bram[2466] = 6'b001000;
frog_bram[2467] = 6'b001100;
frog_bram[2468] = 6'b001100;
frog_bram[2469] = 6'b001100;
frog_bram[2470] = 6'b001100;
frog_bram[2471] = 6'b110000;
frog_bram[2472] = 6'b110000;
frog_bram[2473] = 6'b001100;
frog_bram[2474] = 6'b001100;
frog_bram[2475] = 6'b001100;
frog_bram[2476] = 6'b001100;
frog_bram[2477] = 6'b001000;
frog_bram[2478] = 6'b001100;
frog_bram[2479] = 6'b001100;
frog_bram[2480] = 6'b001100;
frog_bram[2481] = 6'b001000;
frog_bram[2482] = 6'b001100;
frog_bram[2483] = 6'b001100;
frog_bram[2484] = 6'b001100;
frog_bram[2485] = 6'b001000;
frog_bram[2486] = 6'b001000;
frog_bram[2487] = 6'b001100;
frog_bram[2488] = 6'b001100;
frog_bram[2489] = 6'b001000;
frog_bram[2490] = 6'b001000;
frog_bram[2491] = 6'b001000;
frog_bram[2492] = 6'b000000;
frog_bram[2493] = 6'b000000;
frog_bram[2494] = 6'b000000;
frog_bram[2495] = 6'b000000;
frog_bram[2496] = 6'b000000;
frog_bram[2497] = 6'b000000;
frog_bram[2498] = 6'b001000;
frog_bram[2499] = 6'b000100;
frog_bram[2500] = 6'b001100;
frog_bram[2501] = 6'b001100;
frog_bram[2502] = 6'b001100;
frog_bram[2503] = 6'b001100;
frog_bram[2504] = 6'b001100;
frog_bram[2505] = 6'b001100;
frog_bram[2506] = 6'b001100;
frog_bram[2507] = 6'b001100;
frog_bram[2508] = 6'b001100;
frog_bram[2509] = 6'b001000;
frog_bram[2510] = 6'b001100;
frog_bram[2511] = 6'b001100;
frog_bram[2512] = 6'b001000;
frog_bram[2513] = 6'b001000;
frog_bram[2514] = 6'b001000;
frog_bram[2515] = 6'b001000;
frog_bram[2516] = 6'b001000;
frog_bram[2517] = 6'b001000;
frog_bram[2518] = 6'b001000;
frog_bram[2519] = 6'b001000;
frog_bram[2520] = 6'b001000;
frog_bram[2521] = 6'b001000;
frog_bram[2522] = 6'b001000;
frog_bram[2523] = 6'b001000;
frog_bram[2524] = 6'b000000;
frog_bram[2525] = 6'b000000;
frog_bram[2526] = 6'b000000;
frog_bram[2527] = 6'b000000;
frog_bram[2528] = 6'b000000;
frog_bram[2529] = 6'b000000;
frog_bram[2530] = 6'b001100;
frog_bram[2531] = 6'b001100;
frog_bram[2532] = 6'b001100;
frog_bram[2533] = 6'b001100;
frog_bram[2534] = 6'b001100;
frog_bram[2535] = 6'b001100;
frog_bram[2536] = 6'b001100;
frog_bram[2537] = 6'b001100;
frog_bram[2538] = 6'b001100;
frog_bram[2539] = 6'b001100;
frog_bram[2540] = 6'b001100;
frog_bram[2541] = 6'b001000;
frog_bram[2542] = 6'b001000;
frog_bram[2543] = 6'b001000;
frog_bram[2544] = 6'b001000;
frog_bram[2545] = 6'b001000;
frog_bram[2546] = 6'b001000;
frog_bram[2547] = 6'b001000;
frog_bram[2548] = 6'b001000;
frog_bram[2549] = 6'b001000;
frog_bram[2550] = 6'b001000;
frog_bram[2551] = 6'b001000;
frog_bram[2552] = 6'b001000;
frog_bram[2553] = 6'b001000;
frog_bram[2554] = 6'b001000;
frog_bram[2555] = 6'b001000;
frog_bram[2556] = 6'b001000;
frog_bram[2557] = 6'b000000;
frog_bram[2558] = 6'b000000;
frog_bram[2559] = 6'b000000;
frog_bram[2560] = 6'b000000;
frog_bram[2561] = 6'b000000;
frog_bram[2562] = 6'b001100;
frog_bram[2563] = 6'b001100;
frog_bram[2564] = 6'b001100;
frog_bram[2565] = 6'b001100;
frog_bram[2566] = 6'b001100;
frog_bram[2567] = 6'b001100;
frog_bram[2568] = 6'b001100;
frog_bram[2569] = 6'b001100;
frog_bram[2570] = 6'b001100;
frog_bram[2571] = 6'b001100;
frog_bram[2572] = 6'b001100;
frog_bram[2573] = 6'b001000;
frog_bram[2574] = 6'b001000;
frog_bram[2575] = 6'b001000;
frog_bram[2576] = 6'b001000;
frog_bram[2577] = 6'b001000;
frog_bram[2578] = 6'b001000;
frog_bram[2579] = 6'b001000;
frog_bram[2580] = 6'b001000;
frog_bram[2581] = 6'b001000;
frog_bram[2582] = 6'b001000;
frog_bram[2583] = 6'b001000;
frog_bram[2584] = 6'b001000;
frog_bram[2585] = 6'b001000;
frog_bram[2586] = 6'b001000;
frog_bram[2587] = 6'b001000;
frog_bram[2588] = 6'b001000;
frog_bram[2589] = 6'b000000;
frog_bram[2590] = 6'b000000;
frog_bram[2591] = 6'b000000;
frog_bram[2592] = 6'b000000;
frog_bram[2593] = 6'b000000;
frog_bram[2594] = 6'b001000;
frog_bram[2595] = 6'b000100;
frog_bram[2596] = 6'b001100;
frog_bram[2597] = 6'b001100;
frog_bram[2598] = 6'b001100;
frog_bram[2599] = 6'b001000;
frog_bram[2600] = 6'b001000;
frog_bram[2601] = 6'b001000;
frog_bram[2602] = 6'b001100;
frog_bram[2603] = 6'b001100;
frog_bram[2604] = 6'b001100;
frog_bram[2605] = 6'b001000;
frog_bram[2606] = 6'b001100;
frog_bram[2607] = 6'b001100;
frog_bram[2608] = 6'b001000;
frog_bram[2609] = 6'b001000;
frog_bram[2610] = 6'b001000;
frog_bram[2611] = 6'b001000;
frog_bram[2612] = 6'b001000;
frog_bram[2613] = 6'b001000;
frog_bram[2614] = 6'b001000;
frog_bram[2615] = 6'b001000;
frog_bram[2616] = 6'b001000;
frog_bram[2617] = 6'b001000;
frog_bram[2618] = 6'b001000;
frog_bram[2619] = 6'b001000;
frog_bram[2620] = 6'b000000;
frog_bram[2621] = 6'b000000;
frog_bram[2622] = 6'b000000;
frog_bram[2623] = 6'b000000;
frog_bram[2624] = 6'b000000;
frog_bram[2625] = 6'b000000;
frog_bram[2626] = 6'b001000;
frog_bram[2627] = 6'b001100;
frog_bram[2628] = 6'b001100;
frog_bram[2629] = 6'b001100;
frog_bram[2630] = 6'b001000;
frog_bram[2631] = 6'b110000;
frog_bram[2632] = 6'b110000;
frog_bram[2633] = 6'b001000;
frog_bram[2634] = 6'b001000;
frog_bram[2635] = 6'b001100;
frog_bram[2636] = 6'b001100;
frog_bram[2637] = 6'b001100;
frog_bram[2638] = 6'b001100;
frog_bram[2639] = 6'b001100;
frog_bram[2640] = 6'b001100;
frog_bram[2641] = 6'b001000;
frog_bram[2642] = 6'b001100;
frog_bram[2643] = 6'b001100;
frog_bram[2644] = 6'b001100;
frog_bram[2645] = 6'b001000;
frog_bram[2646] = 6'b001000;
frog_bram[2647] = 6'b001100;
frog_bram[2648] = 6'b001100;
frog_bram[2649] = 6'b001000;
frog_bram[2650] = 6'b001000;
frog_bram[2651] = 6'b001000;
frog_bram[2652] = 6'b000000;
frog_bram[2653] = 6'b000000;
frog_bram[2654] = 6'b000000;
frog_bram[2655] = 6'b000000;
frog_bram[2656] = 6'b000000;
frog_bram[2657] = 6'b000000;
frog_bram[2658] = 6'b000000;
frog_bram[2659] = 6'b001100;
frog_bram[2660] = 6'b001100;
frog_bram[2661] = 6'b001000;
frog_bram[2662] = 6'b110000;
frog_bram[2663] = 6'b010000;
frog_bram[2664] = 6'b010000;
frog_bram[2665] = 6'b110000;
frog_bram[2666] = 6'b001000;
frog_bram[2667] = 6'b001100;
frog_bram[2668] = 6'b001100;
frog_bram[2669] = 6'b001100;
frog_bram[2670] = 6'b001100;
frog_bram[2671] = 6'b001100;
frog_bram[2672] = 6'b001100;
frog_bram[2673] = 6'b001100;
frog_bram[2674] = 6'b001100;
frog_bram[2675] = 6'b001100;
frog_bram[2676] = 6'b001100;
frog_bram[2677] = 6'b001000;
frog_bram[2678] = 6'b001000;
frog_bram[2679] = 6'b001100;
frog_bram[2680] = 6'b001100;
frog_bram[2681] = 6'b001100;
frog_bram[2682] = 6'b001000;
frog_bram[2683] = 6'b000000;
frog_bram[2684] = 6'b000000;
frog_bram[2685] = 6'b000000;
frog_bram[2686] = 6'b000000;
frog_bram[2687] = 6'b000000;
frog_bram[2688] = 6'b000000;
frog_bram[2689] = 6'b000000;
frog_bram[2690] = 6'b000000;
frog_bram[2691] = 6'b000000;
frog_bram[2692] = 6'b001000;
frog_bram[2693] = 6'b001000;
frog_bram[2694] = 6'b110000;
frog_bram[2695] = 6'b010000;
frog_bram[2696] = 6'b010000;
frog_bram[2697] = 6'b110000;
frog_bram[2698] = 6'b001000;
frog_bram[2699] = 6'b001100;
frog_bram[2700] = 6'b001100;
frog_bram[2701] = 6'b001100;
frog_bram[2702] = 6'b001100;
frog_bram[2703] = 6'b001100;
frog_bram[2704] = 6'b001100;
frog_bram[2705] = 6'b001100;
frog_bram[2706] = 6'b001100;
frog_bram[2707] = 6'b001100;
frog_bram[2708] = 6'b001100;
frog_bram[2709] = 6'b001100;
frog_bram[2710] = 6'b001000;
frog_bram[2711] = 6'b001100;
frog_bram[2712] = 6'b001100;
frog_bram[2713] = 6'b001000;
frog_bram[2714] = 6'b001000;
frog_bram[2715] = 6'b000000;
frog_bram[2716] = 6'b000000;
frog_bram[2717] = 6'b000000;
frog_bram[2718] = 6'b000000;
frog_bram[2719] = 6'b000000;
frog_bram[2720] = 6'b000000;
frog_bram[2721] = 6'b000000;
frog_bram[2722] = 6'b000000;
frog_bram[2723] = 6'b000000;
frog_bram[2724] = 6'b000000;
frog_bram[2725] = 6'b001000;
frog_bram[2726] = 6'b001000;
frog_bram[2727] = 6'b110000;
frog_bram[2728] = 6'b100000;
frog_bram[2729] = 6'b001000;
frog_bram[2730] = 6'b001100;
frog_bram[2731] = 6'b001100;
frog_bram[2732] = 6'b001000;
frog_bram[2733] = 6'b001000;
frog_bram[2734] = 6'b001100;
frog_bram[2735] = 6'b001100;
frog_bram[2736] = 6'b001100;
frog_bram[2737] = 6'b001100;
frog_bram[2738] = 6'b001100;
frog_bram[2739] = 6'b001100;
frog_bram[2740] = 6'b001100;
frog_bram[2741] = 6'b001100;
frog_bram[2742] = 6'b001000;
frog_bram[2743] = 6'b001000;
frog_bram[2744] = 6'b001000;
frog_bram[2745] = 6'b000000;
frog_bram[2746] = 6'b000000;
frog_bram[2747] = 6'b000000;
frog_bram[2748] = 6'b000000;
frog_bram[2749] = 6'b000000;
frog_bram[2750] = 6'b000000;
frog_bram[2751] = 6'b000000;
frog_bram[2752] = 6'b000000;
frog_bram[2753] = 6'b000000;
frog_bram[2754] = 6'b000000;
frog_bram[2755] = 6'b000000;
frog_bram[2756] = 6'b000000;
frog_bram[2757] = 6'b000000;
frog_bram[2758] = 6'b001000;
frog_bram[2759] = 6'b001000;
frog_bram[2760] = 6'b001000;
frog_bram[2761] = 6'b001100;
frog_bram[2762] = 6'b001100;
frog_bram[2763] = 6'b001100;
frog_bram[2764] = 6'b000000;
frog_bram[2765] = 6'b000000;
frog_bram[2766] = 6'b001000;
frog_bram[2767] = 6'b001100;
frog_bram[2768] = 6'b001100;
frog_bram[2769] = 6'b001100;
frog_bram[2770] = 6'b001100;
frog_bram[2771] = 6'b001100;
frog_bram[2772] = 6'b001000;
frog_bram[2773] = 6'b001000;
frog_bram[2774] = 6'b000000;
frog_bram[2775] = 6'b000000;
frog_bram[2776] = 6'b000000;
frog_bram[2777] = 6'b001000;
frog_bram[2778] = 6'b001000;
frog_bram[2779] = 6'b001000;
frog_bram[2780] = 6'b000000;
frog_bram[2781] = 6'b000000;
frog_bram[2782] = 6'b000000;
frog_bram[2783] = 6'b000000;
frog_bram[2784] = 6'b000000;
frog_bram[2785] = 6'b000000;
frog_bram[2786] = 6'b000000;
frog_bram[2787] = 6'b000000;
frog_bram[2788] = 6'b000000;
frog_bram[2789] = 6'b000000;
frog_bram[2790] = 6'b000000;
frog_bram[2791] = 6'b000000;
frog_bram[2792] = 6'b001000;
frog_bram[2793] = 6'b001100;
frog_bram[2794] = 6'b001100;
frog_bram[2795] = 6'b000000;
frog_bram[2796] = 6'b000000;
frog_bram[2797] = 6'b001000;
frog_bram[2798] = 6'b001100;
frog_bram[2799] = 6'b000000;
frog_bram[2800] = 6'b000000;
frog_bram[2801] = 6'b001000;
frog_bram[2802] = 6'b000000;
frog_bram[2803] = 6'b000000;
frog_bram[2804] = 6'b000000;
frog_bram[2805] = 6'b000000;
frog_bram[2806] = 6'b001000;
frog_bram[2807] = 6'b001000;
frog_bram[2808] = 6'b001000;
frog_bram[2809] = 6'b001100;
frog_bram[2810] = 6'b001100;
frog_bram[2811] = 6'b001100;
frog_bram[2812] = 6'b001100;
frog_bram[2813] = 6'b001000;
frog_bram[2814] = 6'b000000;
frog_bram[2815] = 6'b000000;
frog_bram[2816] = 6'b000000;
frog_bram[2817] = 6'b000000;
frog_bram[2818] = 6'b000000;
frog_bram[2819] = 6'b001000;
frog_bram[2820] = 6'b001000;
frog_bram[2821] = 6'b000000;
frog_bram[2822] = 6'b000000;
frog_bram[2823] = 6'b000000;
frog_bram[2824] = 6'b000000;
frog_bram[2825] = 6'b000000;
frog_bram[2826] = 6'b000000;
frog_bram[2827] = 6'b000000;
frog_bram[2828] = 6'b001000;
frog_bram[2829] = 6'b001000;
frog_bram[2830] = 6'b001000;
frog_bram[2831] = 6'b001100;
frog_bram[2832] = 6'b001000;
frog_bram[2833] = 6'b000000;
frog_bram[2834] = 6'b001000;
frog_bram[2835] = 6'b001000;
frog_bram[2836] = 6'b001000;
frog_bram[2837] = 6'b001000;
frog_bram[2838] = 6'b001100;
frog_bram[2839] = 6'b001100;
frog_bram[2840] = 6'b001100;
frog_bram[2841] = 6'b001100;
frog_bram[2842] = 6'b001100;
frog_bram[2843] = 6'b001100;
frog_bram[2844] = 6'b001100;
frog_bram[2845] = 6'b001100;
frog_bram[2846] = 6'b000000;
frog_bram[2847] = 6'b000000;
frog_bram[2848] = 6'b000000;
frog_bram[2849] = 6'b000000;
frog_bram[2850] = 6'b000000;
frog_bram[2851] = 6'b001000;
frog_bram[2852] = 6'b001100;
frog_bram[2853] = 6'b001100;
frog_bram[2854] = 6'b000000;
frog_bram[2855] = 6'b001000;
frog_bram[2856] = 6'b001000;
frog_bram[2857] = 6'b000000;
frog_bram[2858] = 6'b000000;
frog_bram[2859] = 6'b000000;
frog_bram[2860] = 6'b001000;
frog_bram[2861] = 6'b001000;
frog_bram[2862] = 6'b001000;
frog_bram[2863] = 6'b001000;
frog_bram[2864] = 6'b000000;
frog_bram[2865] = 6'b000000;
frog_bram[2866] = 6'b001000;
frog_bram[2867] = 6'b001100;
frog_bram[2868] = 6'b001100;
frog_bram[2869] = 6'b001100;
frog_bram[2870] = 6'b001100;
frog_bram[2871] = 6'b001100;
frog_bram[2872] = 6'b001000;
frog_bram[2873] = 6'b001000;
frog_bram[2874] = 6'b000000;
frog_bram[2875] = 6'b001100;
frog_bram[2876] = 6'b001100;
frog_bram[2877] = 6'b001100;
frog_bram[2878] = 6'b001000;
frog_bram[2879] = 6'b000000;
frog_bram[2880] = 6'b000000;
frog_bram[2881] = 6'b000000;
frog_bram[2882] = 6'b000000;
frog_bram[2883] = 6'b000000;
frog_bram[2884] = 6'b000000;
frog_bram[2885] = 6'b001100;
frog_bram[2886] = 6'b001000;
frog_bram[2887] = 6'b000100;
frog_bram[2888] = 6'b001100;
frog_bram[2889] = 6'b001100;
frog_bram[2890] = 6'b000000;
frog_bram[2891] = 6'b001000;
frog_bram[2892] = 6'b001000;
frog_bram[2893] = 6'b001000;
frog_bram[2894] = 6'b001000;
frog_bram[2895] = 6'b000000;
frog_bram[2896] = 6'b000000;
frog_bram[2897] = 6'b000000;
frog_bram[2898] = 6'b000000;
frog_bram[2899] = 6'b001000;
frog_bram[2900] = 6'b001000;
frog_bram[2901] = 6'b001000;
frog_bram[2902] = 6'b001000;
frog_bram[2903] = 6'b001000;
frog_bram[2904] = 6'b001000;
frog_bram[2905] = 6'b000000;
frog_bram[2906] = 6'b001000;
frog_bram[2907] = 6'b001100;
frog_bram[2908] = 6'b001100;
frog_bram[2909] = 6'b001100;
frog_bram[2910] = 6'b001000;
frog_bram[2911] = 6'b000000;
frog_bram[2912] = 6'b000000;
frog_bram[2913] = 6'b000000;
frog_bram[2914] = 6'b000000;
frog_bram[2915] = 6'b001000;
frog_bram[2916] = 6'b001000;
frog_bram[2917] = 6'b000100;
frog_bram[2918] = 6'b001000;
frog_bram[2919] = 6'b001100;
frog_bram[2920] = 6'b001100;
frog_bram[2921] = 6'b001100;
frog_bram[2922] = 6'b001100;
frog_bram[2923] = 6'b001100;
frog_bram[2924] = 6'b001100;
frog_bram[2925] = 6'b001000;
frog_bram[2926] = 6'b001000;
frog_bram[2927] = 6'b000000;
frog_bram[2928] = 6'b000000;
frog_bram[2929] = 6'b000000;
frog_bram[2930] = 6'b000000;
frog_bram[2931] = 6'b000000;
frog_bram[2932] = 6'b000000;
frog_bram[2933] = 6'b000000;
frog_bram[2934] = 6'b000000;
frog_bram[2935] = 6'b000000;
frog_bram[2936] = 6'b000000;
frog_bram[2937] = 6'b001000;
frog_bram[2938] = 6'b001100;
frog_bram[2939] = 6'b001100;
frog_bram[2940] = 6'b001100;
frog_bram[2941] = 6'b001000;
frog_bram[2942] = 6'b000000;
frog_bram[2943] = 6'b000000;
frog_bram[2944] = 6'b000000;
frog_bram[2945] = 6'b000000;
frog_bram[2946] = 6'b000000;
frog_bram[2947] = 6'b001100;
frog_bram[2948] = 6'b001100;
frog_bram[2949] = 6'b001100;
frog_bram[2950] = 6'b001100;
frog_bram[2951] = 6'b001100;
frog_bram[2952] = 6'b001100;
frog_bram[2953] = 6'b001100;
frog_bram[2954] = 6'b001100;
frog_bram[2955] = 6'b001100;
frog_bram[2956] = 6'b001100;
frog_bram[2957] = 6'b001000;
frog_bram[2958] = 6'b000000;
frog_bram[2959] = 6'b000000;
frog_bram[2960] = 6'b000000;
frog_bram[2961] = 6'b000000;
frog_bram[2962] = 6'b000000;
frog_bram[2963] = 6'b000000;
frog_bram[2964] = 6'b000000;
frog_bram[2965] = 6'b000000;
frog_bram[2966] = 6'b001000;
frog_bram[2967] = 6'b001100;
frog_bram[2968] = 6'b001100;
frog_bram[2969] = 6'b001100;
frog_bram[2970] = 6'b001100;
frog_bram[2971] = 6'b001100;
frog_bram[2972] = 6'b001100;
frog_bram[2973] = 6'b001000;
frog_bram[2974] = 6'b000000;
frog_bram[2975] = 6'b000000;
frog_bram[2976] = 6'b000000;
frog_bram[2977] = 6'b000000;
frog_bram[2978] = 6'b000000;
frog_bram[2979] = 6'b000000;
frog_bram[2980] = 6'b000000;
frog_bram[2981] = 6'b000000;
frog_bram[2982] = 6'b000000;
frog_bram[2983] = 6'b001100;
frog_bram[2984] = 6'b001100;
frog_bram[2985] = 6'b001100;
frog_bram[2986] = 6'b001100;
frog_bram[2987] = 6'b001100;
frog_bram[2988] = 6'b001100;
frog_bram[2989] = 6'b000000;
frog_bram[2990] = 6'b000000;
frog_bram[2991] = 6'b000000;
frog_bram[2992] = 6'b000000;
frog_bram[2993] = 6'b000000;
frog_bram[2994] = 6'b000000;
frog_bram[2995] = 6'b000000;
frog_bram[2996] = 6'b000000;
frog_bram[2997] = 6'b000000;
frog_bram[2998] = 6'b001000;
frog_bram[2999] = 6'b001100;
frog_bram[3000] = 6'b000100;
frog_bram[3001] = 6'b001000;
frog_bram[3002] = 6'b001100;
frog_bram[3003] = 6'b001100;
frog_bram[3004] = 6'b001100;
frog_bram[3005] = 6'b001000;
frog_bram[3006] = 6'b000000;
frog_bram[3007] = 6'b000000;
frog_bram[3008] = 6'b000000;
frog_bram[3009] = 6'b000000;
frog_bram[3010] = 6'b000000;
frog_bram[3011] = 6'b000000;
frog_bram[3012] = 6'b000000;
frog_bram[3013] = 6'b000000;
frog_bram[3014] = 6'b000000;
frog_bram[3015] = 6'b000000;
frog_bram[3016] = 6'b000000;
frog_bram[3017] = 6'b000000;
frog_bram[3018] = 6'b000000;
frog_bram[3019] = 6'b000000;
frog_bram[3020] = 6'b000000;
frog_bram[3021] = 6'b000000;
frog_bram[3022] = 6'b000000;
frog_bram[3023] = 6'b000000;
frog_bram[3024] = 6'b000000;
frog_bram[3025] = 6'b000000;
frog_bram[3026] = 6'b000000;
frog_bram[3027] = 6'b000000;
frog_bram[3028] = 6'b000000;
frog_bram[3029] = 6'b000000;
frog_bram[3030] = 6'b000000;
frog_bram[3031] = 6'b000000;
frog_bram[3032] = 6'b001000;
frog_bram[3033] = 6'b001100;
frog_bram[3034] = 6'b001100;
frog_bram[3035] = 6'b001100;
frog_bram[3036] = 6'b001100;
frog_bram[3037] = 6'b000000;
frog_bram[3038] = 6'b000000;
frog_bram[3039] = 6'b000000;
frog_bram[3040] = 6'b000000;
frog_bram[3041] = 6'b000000;
frog_bram[3042] = 6'b000000;
frog_bram[3043] = 6'b000000;
frog_bram[3044] = 6'b000000;
frog_bram[3045] = 6'b000000;
frog_bram[3046] = 6'b000000;
frog_bram[3047] = 6'b000000;
frog_bram[3048] = 6'b000000;
frog_bram[3049] = 6'b000000;
frog_bram[3050] = 6'b000000;
frog_bram[3051] = 6'b000000;
frog_bram[3052] = 6'b000000;
frog_bram[3053] = 6'b000000;
frog_bram[3054] = 6'b000000;
frog_bram[3055] = 6'b000000;
frog_bram[3056] = 6'b000000;
frog_bram[3057] = 6'b000000;
frog_bram[3058] = 6'b000000;
frog_bram[3059] = 6'b000000;
frog_bram[3060] = 6'b000000;
frog_bram[3061] = 6'b000000;
frog_bram[3062] = 6'b000000;
frog_bram[3063] = 6'b000000;
frog_bram[3064] = 6'b001000;
frog_bram[3065] = 6'b001100;
frog_bram[3066] = 6'b000000;
frog_bram[3067] = 6'b001000;
frog_bram[3068] = 6'b001100;
frog_bram[3069] = 6'b000000;
frog_bram[3070] = 6'b000000;
frog_bram[3071] = 6'b000000;
        // Add more initialization here for the right-facing sprite (3072 - 4095)
frog_bram[3072] = 6'b000000;
frog_bram[3073] = 6'b000000;
frog_bram[3074] = 6'b000000;
frog_bram[3075] = 6'b001100;
frog_bram[3076] = 6'b001000;
frog_bram[3077] = 6'b000000;
frog_bram[3078] = 6'b001100;
frog_bram[3079] = 6'b001000;
frog_bram[3080] = 6'b000000;
frog_bram[3081] = 6'b000000;
frog_bram[3082] = 6'b000000;
frog_bram[3083] = 6'b000000;
frog_bram[3084] = 6'b000000;
frog_bram[3085] = 6'b000000;
frog_bram[3086] = 6'b000000;
frog_bram[3087] = 6'b000000;
frog_bram[3088] = 6'b000000;
frog_bram[3089] = 6'b000000;
frog_bram[3090] = 6'b000000;
frog_bram[3091] = 6'b000000;
frog_bram[3092] = 6'b000000;
frog_bram[3093] = 6'b000000;
frog_bram[3094] = 6'b000000;
frog_bram[3095] = 6'b000000;
frog_bram[3096] = 6'b000000;
frog_bram[3097] = 6'b000000;
frog_bram[3098] = 6'b000000;
frog_bram[3099] = 6'b000000;
frog_bram[3100] = 6'b000000;
frog_bram[3101] = 6'b000000;
frog_bram[3102] = 6'b000000;
frog_bram[3103] = 6'b000000;
frog_bram[3104] = 6'b000000;
frog_bram[3105] = 6'b000000;
frog_bram[3106] = 6'b000000;
frog_bram[3107] = 6'b001100;
frog_bram[3108] = 6'b001100;
frog_bram[3109] = 6'b001100;
frog_bram[3110] = 6'b001100;
frog_bram[3111] = 6'b001000;
frog_bram[3112] = 6'b000000;
frog_bram[3113] = 6'b000000;
frog_bram[3114] = 6'b000000;
frog_bram[3115] = 6'b000000;
frog_bram[3116] = 6'b000000;
frog_bram[3117] = 6'b000000;
frog_bram[3118] = 6'b000000;
frog_bram[3119] = 6'b000000;
frog_bram[3120] = 6'b000000;
frog_bram[3121] = 6'b000000;
frog_bram[3122] = 6'b000000;
frog_bram[3123] = 6'b000000;
frog_bram[3124] = 6'b000000;
frog_bram[3125] = 6'b000000;
frog_bram[3126] = 6'b000000;
frog_bram[3127] = 6'b000000;
frog_bram[3128] = 6'b000000;
frog_bram[3129] = 6'b000000;
frog_bram[3130] = 6'b000000;
frog_bram[3131] = 6'b000000;
frog_bram[3132] = 6'b000000;
frog_bram[3133] = 6'b000000;
frog_bram[3134] = 6'b000000;
frog_bram[3135] = 6'b000000;
frog_bram[3136] = 6'b000000;
frog_bram[3137] = 6'b000000;
frog_bram[3138] = 6'b001000;
frog_bram[3139] = 6'b001100;
frog_bram[3140] = 6'b001100;
frog_bram[3141] = 6'b001100;
frog_bram[3142] = 6'b001000;
frog_bram[3143] = 6'b000100;
frog_bram[3144] = 6'b001100;
frog_bram[3145] = 6'b001000;
frog_bram[3146] = 6'b000000;
frog_bram[3147] = 6'b000000;
frog_bram[3148] = 6'b000000;
frog_bram[3149] = 6'b000000;
frog_bram[3150] = 6'b000000;
frog_bram[3151] = 6'b000000;
frog_bram[3152] = 6'b000000;
frog_bram[3153] = 6'b000000;
frog_bram[3154] = 6'b000000;
frog_bram[3155] = 6'b001100;
frog_bram[3156] = 6'b001100;
frog_bram[3157] = 6'b001100;
frog_bram[3158] = 6'b001100;
frog_bram[3159] = 6'b001100;
frog_bram[3160] = 6'b001100;
frog_bram[3161] = 6'b000000;
frog_bram[3162] = 6'b000000;
frog_bram[3163] = 6'b000000;
frog_bram[3164] = 6'b000000;
frog_bram[3165] = 6'b000000;
frog_bram[3166] = 6'b000000;
frog_bram[3167] = 6'b000000;
frog_bram[3168] = 6'b000000;
frog_bram[3169] = 6'b000000;
frog_bram[3170] = 6'b001000;
frog_bram[3171] = 6'b001100;
frog_bram[3172] = 6'b001100;
frog_bram[3173] = 6'b001100;
frog_bram[3174] = 6'b001100;
frog_bram[3175] = 6'b001100;
frog_bram[3176] = 6'b001100;
frog_bram[3177] = 6'b001000;
frog_bram[3178] = 6'b000000;
frog_bram[3179] = 6'b000000;
frog_bram[3180] = 6'b000000;
frog_bram[3181] = 6'b000000;
frog_bram[3182] = 6'b000000;
frog_bram[3183] = 6'b000000;
frog_bram[3184] = 6'b000000;
frog_bram[3185] = 6'b000000;
frog_bram[3186] = 6'b001000;
frog_bram[3187] = 6'b001100;
frog_bram[3188] = 6'b001100;
frog_bram[3189] = 6'b001100;
frog_bram[3190] = 6'b001100;
frog_bram[3191] = 6'b001100;
frog_bram[3192] = 6'b001100;
frog_bram[3193] = 6'b001100;
frog_bram[3194] = 6'b001100;
frog_bram[3195] = 6'b001100;
frog_bram[3196] = 6'b001100;
frog_bram[3197] = 6'b000000;
frog_bram[3198] = 6'b000000;
frog_bram[3199] = 6'b000000;
frog_bram[3200] = 6'b000000;
frog_bram[3201] = 6'b000000;
frog_bram[3202] = 6'b001000;
frog_bram[3203] = 6'b001100;
frog_bram[3204] = 6'b001100;
frog_bram[3205] = 6'b001100;
frog_bram[3206] = 6'b001000;
frog_bram[3207] = 6'b000000;
frog_bram[3208] = 6'b000000;
frog_bram[3209] = 6'b000000;
frog_bram[3210] = 6'b000000;
frog_bram[3211] = 6'b000000;
frog_bram[3212] = 6'b000000;
frog_bram[3213] = 6'b000000;
frog_bram[3214] = 6'b000000;
frog_bram[3215] = 6'b000000;
frog_bram[3216] = 6'b000000;
frog_bram[3217] = 6'b001000;
frog_bram[3218] = 6'b001000;
frog_bram[3219] = 6'b001100;
frog_bram[3220] = 6'b001100;
frog_bram[3221] = 6'b001100;
frog_bram[3222] = 6'b001100;
frog_bram[3223] = 6'b001100;
frog_bram[3224] = 6'b001100;
frog_bram[3225] = 6'b001000;
frog_bram[3226] = 6'b000100;
frog_bram[3227] = 6'b001000;
frog_bram[3228] = 6'b001000;
frog_bram[3229] = 6'b000000;
frog_bram[3230] = 6'b000000;
frog_bram[3231] = 6'b000000;
frog_bram[3232] = 6'b000000;
frog_bram[3233] = 6'b001000;
frog_bram[3234] = 6'b001100;
frog_bram[3235] = 6'b001100;
frog_bram[3236] = 6'b001100;
frog_bram[3237] = 6'b001000;
frog_bram[3238] = 6'b000000;
frog_bram[3239] = 6'b001000;
frog_bram[3240] = 6'b001000;
frog_bram[3241] = 6'b001000;
frog_bram[3242] = 6'b001000;
frog_bram[3243] = 6'b001000;
frog_bram[3244] = 6'b001000;
frog_bram[3245] = 6'b000000;
frog_bram[3246] = 6'b000000;
frog_bram[3247] = 6'b000000;
frog_bram[3248] = 6'b000000;
frog_bram[3249] = 6'b001000;
frog_bram[3250] = 6'b001000;
frog_bram[3251] = 6'b001000;
frog_bram[3252] = 6'b001000;
frog_bram[3253] = 6'b000000;
frog_bram[3254] = 6'b001100;
frog_bram[3255] = 6'b001100;
frog_bram[3256] = 6'b000100;
frog_bram[3257] = 6'b001000;
frog_bram[3258] = 6'b001100;
frog_bram[3259] = 6'b000000;
frog_bram[3260] = 6'b000000;
frog_bram[3261] = 6'b000000;
frog_bram[3262] = 6'b000000;
frog_bram[3263] = 6'b000000;
frog_bram[3264] = 6'b000000;
frog_bram[3265] = 6'b001000;
frog_bram[3266] = 6'b001100;
frog_bram[3267] = 6'b001100;
frog_bram[3268] = 6'b001100;
frog_bram[3269] = 6'b000000;
frog_bram[3270] = 6'b001000;
frog_bram[3271] = 6'b001000;
frog_bram[3272] = 6'b001100;
frog_bram[3273] = 6'b001100;
frog_bram[3274] = 6'b001100;
frog_bram[3275] = 6'b001100;
frog_bram[3276] = 6'b001100;
frog_bram[3277] = 6'b001000;
frog_bram[3278] = 6'b000000;
frog_bram[3279] = 6'b000000;
frog_bram[3280] = 6'b001000;
frog_bram[3281] = 6'b001000;
frog_bram[3282] = 6'b001000;
frog_bram[3283] = 6'b001000;
frog_bram[3284] = 6'b000000;
frog_bram[3285] = 6'b000000;
frog_bram[3286] = 6'b000000;
frog_bram[3287] = 6'b001000;
frog_bram[3288] = 6'b001000;
frog_bram[3289] = 6'b000000;
frog_bram[3290] = 6'b001100;
frog_bram[3291] = 6'b001100;
frog_bram[3292] = 6'b001000;
frog_bram[3293] = 6'b000000;
frog_bram[3294] = 6'b000000;
frog_bram[3295] = 6'b000000;
frog_bram[3296] = 6'b000000;
frog_bram[3297] = 6'b000000;
frog_bram[3298] = 6'b001100;
frog_bram[3299] = 6'b001100;
frog_bram[3300] = 6'b001100;
frog_bram[3301] = 6'b001100;
frog_bram[3302] = 6'b001100;
frog_bram[3303] = 6'b001100;
frog_bram[3304] = 6'b001100;
frog_bram[3305] = 6'b001100;
frog_bram[3306] = 6'b001000;
frog_bram[3307] = 6'b001000;
frog_bram[3308] = 6'b001000;
frog_bram[3309] = 6'b001000;
frog_bram[3310] = 6'b000000;
frog_bram[3311] = 6'b001000;
frog_bram[3312] = 6'b001100;
frog_bram[3313] = 6'b001000;
frog_bram[3314] = 6'b001000;
frog_bram[3315] = 6'b001000;
frog_bram[3316] = 6'b000000;
frog_bram[3317] = 6'b000000;
frog_bram[3318] = 6'b000000;
frog_bram[3319] = 6'b000000;
frog_bram[3320] = 6'b000000;
frog_bram[3321] = 6'b000000;
frog_bram[3322] = 6'b000000;
frog_bram[3323] = 6'b001000;
frog_bram[3324] = 6'b001000;
frog_bram[3325] = 6'b000000;
frog_bram[3326] = 6'b000000;
frog_bram[3327] = 6'b000000;
frog_bram[3328] = 6'b000000;
frog_bram[3329] = 6'b000000;
frog_bram[3330] = 6'b001000;
frog_bram[3331] = 6'b001100;
frog_bram[3332] = 6'b001100;
frog_bram[3333] = 6'b001100;
frog_bram[3334] = 6'b001100;
frog_bram[3335] = 6'b001000;
frog_bram[3336] = 6'b001000;
frog_bram[3337] = 6'b001000;
frog_bram[3338] = 6'b000000;
frog_bram[3339] = 6'b000000;
frog_bram[3340] = 6'b000000;
frog_bram[3341] = 6'b000000;
frog_bram[3342] = 6'b001000;
frog_bram[3343] = 6'b000000;
frog_bram[3344] = 6'b000000;
frog_bram[3345] = 6'b001100;
frog_bram[3346] = 6'b001000;
frog_bram[3347] = 6'b000000;
frog_bram[3348] = 6'b000000;
frog_bram[3349] = 6'b001100;
frog_bram[3350] = 6'b001100;
frog_bram[3351] = 6'b001000;
frog_bram[3352] = 6'b000000;
frog_bram[3353] = 6'b000000;
frog_bram[3354] = 6'b000000;
frog_bram[3355] = 6'b000000;
frog_bram[3356] = 6'b000000;
frog_bram[3357] = 6'b000000;
frog_bram[3358] = 6'b000000;
frog_bram[3359] = 6'b000000;
frog_bram[3360] = 6'b000000;
frog_bram[3361] = 6'b000000;
frog_bram[3362] = 6'b000000;
frog_bram[3363] = 6'b000000;
frog_bram[3364] = 6'b001000;
frog_bram[3365] = 6'b001000;
frog_bram[3366] = 6'b001000;
frog_bram[3367] = 6'b000000;
frog_bram[3368] = 6'b000000;
frog_bram[3369] = 6'b000000;
frog_bram[3370] = 6'b001000;
frog_bram[3371] = 6'b001000;
frog_bram[3372] = 6'b001100;
frog_bram[3373] = 6'b001100;
frog_bram[3374] = 6'b001100;
frog_bram[3375] = 6'b001100;
frog_bram[3376] = 6'b001100;
frog_bram[3377] = 6'b001000;
frog_bram[3378] = 6'b000000;
frog_bram[3379] = 6'b000000;
frog_bram[3380] = 6'b001100;
frog_bram[3381] = 6'b001100;
frog_bram[3382] = 6'b001100;
frog_bram[3383] = 6'b001000;
frog_bram[3384] = 6'b001000;
frog_bram[3385] = 6'b001000;
frog_bram[3386] = 6'b000000;
frog_bram[3387] = 6'b000000;
frog_bram[3388] = 6'b000000;
frog_bram[3389] = 6'b000000;
frog_bram[3390] = 6'b000000;
frog_bram[3391] = 6'b000000;
frog_bram[3392] = 6'b000000;
frog_bram[3393] = 6'b000000;
frog_bram[3394] = 6'b000000;
frog_bram[3395] = 6'b000000;
frog_bram[3396] = 6'b000000;
frog_bram[3397] = 6'b000000;
frog_bram[3398] = 6'b000000;
frog_bram[3399] = 6'b001000;
frog_bram[3400] = 6'b001000;
frog_bram[3401] = 6'b001000;
frog_bram[3402] = 6'b001100;
frog_bram[3403] = 6'b001100;
frog_bram[3404] = 6'b001100;
frog_bram[3405] = 6'b001100;
frog_bram[3406] = 6'b001100;
frog_bram[3407] = 6'b001100;
frog_bram[3408] = 6'b001100;
frog_bram[3409] = 6'b001100;
frog_bram[3410] = 6'b001000;
frog_bram[3411] = 6'b001000;
frog_bram[3412] = 6'b001100;
frog_bram[3413] = 6'b001100;
frog_bram[3414] = 6'b001000;
frog_bram[3415] = 6'b100000;
frog_bram[3416] = 6'b110000;
frog_bram[3417] = 6'b001000;
frog_bram[3418] = 6'b001000;
frog_bram[3419] = 6'b000000;
frog_bram[3420] = 6'b000000;
frog_bram[3421] = 6'b000000;
frog_bram[3422] = 6'b000000;
frog_bram[3423] = 6'b000000;
frog_bram[3424] = 6'b000000;
frog_bram[3425] = 6'b000000;
frog_bram[3426] = 6'b000000;
frog_bram[3427] = 6'b000000;
frog_bram[3428] = 6'b000000;
frog_bram[3429] = 6'b001000;
frog_bram[3430] = 6'b001000;
frog_bram[3431] = 6'b001100;
frog_bram[3432] = 6'b001100;
frog_bram[3433] = 6'b001000;
frog_bram[3434] = 6'b001100;
frog_bram[3435] = 6'b001100;
frog_bram[3436] = 6'b001100;
frog_bram[3437] = 6'b001100;
frog_bram[3438] = 6'b001100;
frog_bram[3439] = 6'b001100;
frog_bram[3440] = 6'b001100;
frog_bram[3441] = 6'b001100;
frog_bram[3442] = 6'b001100;
frog_bram[3443] = 6'b001100;
frog_bram[3444] = 6'b001100;
frog_bram[3445] = 6'b001000;
frog_bram[3446] = 6'b110000;
frog_bram[3447] = 6'b010000;
frog_bram[3448] = 6'b010000;
frog_bram[3449] = 6'b110000;
frog_bram[3450] = 6'b001000;
frog_bram[3451] = 6'b001000;
frog_bram[3452] = 6'b000000;
frog_bram[3453] = 6'b000000;
frog_bram[3454] = 6'b000000;
frog_bram[3455] = 6'b000000;
frog_bram[3456] = 6'b000000;
frog_bram[3457] = 6'b000000;
frog_bram[3458] = 6'b000000;
frog_bram[3459] = 6'b000000;
frog_bram[3460] = 6'b000000;
frog_bram[3461] = 6'b001000;
frog_bram[3462] = 6'b001100;
frog_bram[3463] = 6'b001100;
frog_bram[3464] = 6'b001100;
frog_bram[3465] = 6'b001000;
frog_bram[3466] = 6'b001000;
frog_bram[3467] = 6'b001100;
frog_bram[3468] = 6'b001100;
frog_bram[3469] = 6'b001100;
frog_bram[3470] = 6'b001100;
frog_bram[3471] = 6'b001100;
frog_bram[3472] = 6'b001100;
frog_bram[3473] = 6'b001100;
frog_bram[3474] = 6'b001100;
frog_bram[3475] = 6'b001100;
frog_bram[3476] = 6'b001100;
frog_bram[3477] = 6'b001000;
frog_bram[3478] = 6'b110000;
frog_bram[3479] = 6'b010000;
frog_bram[3480] = 6'b010000;
frog_bram[3481] = 6'b110000;
frog_bram[3482] = 6'b001000;
frog_bram[3483] = 6'b001100;
frog_bram[3484] = 6'b001100;
frog_bram[3485] = 6'b000000;
frog_bram[3486] = 6'b000000;
frog_bram[3487] = 6'b000000;
frog_bram[3488] = 6'b000000;
frog_bram[3489] = 6'b000000;
frog_bram[3490] = 6'b000000;
frog_bram[3491] = 6'b000000;
frog_bram[3492] = 6'b001000;
frog_bram[3493] = 6'b001000;
frog_bram[3494] = 6'b001000;
frog_bram[3495] = 6'b001100;
frog_bram[3496] = 6'b001100;
frog_bram[3497] = 6'b001000;
frog_bram[3498] = 6'b001000;
frog_bram[3499] = 6'b001100;
frog_bram[3500] = 6'b001100;
frog_bram[3501] = 6'b001100;
frog_bram[3502] = 6'b001000;
frog_bram[3503] = 6'b001100;
frog_bram[3504] = 6'b001100;
frog_bram[3505] = 6'b001100;
frog_bram[3506] = 6'b001100;
frog_bram[3507] = 6'b001100;
frog_bram[3508] = 6'b001100;
frog_bram[3509] = 6'b001000;
frog_bram[3510] = 6'b001000;
frog_bram[3511] = 6'b110000;
frog_bram[3512] = 6'b110000;
frog_bram[3513] = 6'b001000;
frog_bram[3514] = 6'b001100;
frog_bram[3515] = 6'b001100;
frog_bram[3516] = 6'b001100;
frog_bram[3517] = 6'b001000;
frog_bram[3518] = 6'b000000;
frog_bram[3519] = 6'b000000;
frog_bram[3520] = 6'b000000;
frog_bram[3521] = 6'b000000;
frog_bram[3522] = 6'b000000;
frog_bram[3523] = 6'b000000;
frog_bram[3524] = 6'b001000;
frog_bram[3525] = 6'b001000;
frog_bram[3526] = 6'b001000;
frog_bram[3527] = 6'b001000;
frog_bram[3528] = 6'b001000;
frog_bram[3529] = 6'b001000;
frog_bram[3530] = 6'b001000;
frog_bram[3531] = 6'b001000;
frog_bram[3532] = 6'b001000;
frog_bram[3533] = 6'b001000;
frog_bram[3534] = 6'b001000;
frog_bram[3535] = 6'b001000;
frog_bram[3536] = 6'b001100;
frog_bram[3537] = 6'b001100;
frog_bram[3538] = 6'b001000;
frog_bram[3539] = 6'b001100;
frog_bram[3540] = 6'b001100;
frog_bram[3541] = 6'b001100;
frog_bram[3542] = 6'b001000;
frog_bram[3543] = 6'b001000;
frog_bram[3544] = 6'b001000;
frog_bram[3545] = 6'b001100;
frog_bram[3546] = 6'b001100;
frog_bram[3547] = 6'b001100;
frog_bram[3548] = 6'b000100;
frog_bram[3549] = 6'b001000;
frog_bram[3550] = 6'b000000;
frog_bram[3551] = 6'b000000;
frog_bram[3552] = 6'b000000;
frog_bram[3553] = 6'b000000;
frog_bram[3554] = 6'b000000;
frog_bram[3555] = 6'b001000;
frog_bram[3556] = 6'b001000;
frog_bram[3557] = 6'b001000;
frog_bram[3558] = 6'b001000;
frog_bram[3559] = 6'b001000;
frog_bram[3560] = 6'b001000;
frog_bram[3561] = 6'b001000;
frog_bram[3562] = 6'b001000;
frog_bram[3563] = 6'b001000;
frog_bram[3564] = 6'b001000;
frog_bram[3565] = 6'b001000;
frog_bram[3566] = 6'b001000;
frog_bram[3567] = 6'b001000;
frog_bram[3568] = 6'b001000;
frog_bram[3569] = 6'b001000;
frog_bram[3570] = 6'b001000;
frog_bram[3571] = 6'b001100;
frog_bram[3572] = 6'b001100;
frog_bram[3573] = 6'b001100;
frog_bram[3574] = 6'b001100;
frog_bram[3575] = 6'b001100;
frog_bram[3576] = 6'b001100;
frog_bram[3577] = 6'b001100;
frog_bram[3578] = 6'b001100;
frog_bram[3579] = 6'b001100;
frog_bram[3580] = 6'b001100;
frog_bram[3581] = 6'b001100;
frog_bram[3582] = 6'b000000;
frog_bram[3583] = 6'b000000;
frog_bram[3584] = 6'b000000;
frog_bram[3585] = 6'b000000;
frog_bram[3586] = 6'b000000;
frog_bram[3587] = 6'b001000;
frog_bram[3588] = 6'b001000;
frog_bram[3589] = 6'b001000;
frog_bram[3590] = 6'b001000;
frog_bram[3591] = 6'b001000;
frog_bram[3592] = 6'b001000;
frog_bram[3593] = 6'b001000;
frog_bram[3594] = 6'b001000;
frog_bram[3595] = 6'b001000;
frog_bram[3596] = 6'b001000;
frog_bram[3597] = 6'b001000;
frog_bram[3598] = 6'b001000;
frog_bram[3599] = 6'b001000;
frog_bram[3600] = 6'b001000;
frog_bram[3601] = 6'b001000;
frog_bram[3602] = 6'b001000;
frog_bram[3603] = 6'b001100;
frog_bram[3604] = 6'b001100;
frog_bram[3605] = 6'b001100;
frog_bram[3606] = 6'b001100;
frog_bram[3607] = 6'b001100;
frog_bram[3608] = 6'b001100;
frog_bram[3609] = 6'b001100;
frog_bram[3610] = 6'b001100;
frog_bram[3611] = 6'b001100;
frog_bram[3612] = 6'b001100;
frog_bram[3613] = 6'b001100;
frog_bram[3614] = 6'b000000;
frog_bram[3615] = 6'b000000;
frog_bram[3616] = 6'b000000;
frog_bram[3617] = 6'b000000;
frog_bram[3618] = 6'b000000;
frog_bram[3619] = 6'b000000;
frog_bram[3620] = 6'b001000;
frog_bram[3621] = 6'b001000;
frog_bram[3622] = 6'b001000;
frog_bram[3623] = 6'b001000;
frog_bram[3624] = 6'b001000;
frog_bram[3625] = 6'b001000;
frog_bram[3626] = 6'b001000;
frog_bram[3627] = 6'b001000;
frog_bram[3628] = 6'b001000;
frog_bram[3629] = 6'b001000;
frog_bram[3630] = 6'b001000;
frog_bram[3631] = 6'b001000;
frog_bram[3632] = 6'b001100;
frog_bram[3633] = 6'b001100;
frog_bram[3634] = 6'b001000;
frog_bram[3635] = 6'b001100;
frog_bram[3636] = 6'b001100;
frog_bram[3637] = 6'b001100;
frog_bram[3638] = 6'b001100;
frog_bram[3639] = 6'b001100;
frog_bram[3640] = 6'b001100;
frog_bram[3641] = 6'b001100;
frog_bram[3642] = 6'b001100;
frog_bram[3643] = 6'b001100;
frog_bram[3644] = 6'b000100;
frog_bram[3645] = 6'b001000;
frog_bram[3646] = 6'b000000;
frog_bram[3647] = 6'b000000;
frog_bram[3648] = 6'b000000;
frog_bram[3649] = 6'b000000;
frog_bram[3650] = 6'b000000;
frog_bram[3651] = 6'b000000;
frog_bram[3652] = 6'b001000;
frog_bram[3653] = 6'b001000;
frog_bram[3654] = 6'b001000;
frog_bram[3655] = 6'b001100;
frog_bram[3656] = 6'b001100;
frog_bram[3657] = 6'b001000;
frog_bram[3658] = 6'b001000;
frog_bram[3659] = 6'b001100;
frog_bram[3660] = 6'b001100;
frog_bram[3661] = 6'b001100;
frog_bram[3662] = 6'b001000;
frog_bram[3663] = 6'b001100;
frog_bram[3664] = 6'b001100;
frog_bram[3665] = 6'b001100;
frog_bram[3666] = 6'b001000;
frog_bram[3667] = 6'b001100;
frog_bram[3668] = 6'b001100;
frog_bram[3669] = 6'b001100;
frog_bram[3670] = 6'b001100;
frog_bram[3671] = 6'b110000;
frog_bram[3672] = 6'b110000;
frog_bram[3673] = 6'b001100;
frog_bram[3674] = 6'b001100;
frog_bram[3675] = 6'b001100;
frog_bram[3676] = 6'b001100;
frog_bram[3677] = 6'b001000;
frog_bram[3678] = 6'b000000;
frog_bram[3679] = 6'b000000;
frog_bram[3680] = 6'b000000;
frog_bram[3681] = 6'b000000;
frog_bram[3682] = 6'b000000;
frog_bram[3683] = 6'b000000;
frog_bram[3684] = 6'b000000;
frog_bram[3685] = 6'b001000;
frog_bram[3686] = 6'b001100;
frog_bram[3687] = 6'b001100;
frog_bram[3688] = 6'b001100;
frog_bram[3689] = 6'b001000;
frog_bram[3690] = 6'b001000;
frog_bram[3691] = 6'b001100;
frog_bram[3692] = 6'b001100;
frog_bram[3693] = 6'b001100;
frog_bram[3694] = 6'b001100;
frog_bram[3695] = 6'b001100;
frog_bram[3696] = 6'b001100;
frog_bram[3697] = 6'b001100;
frog_bram[3698] = 6'b001100;
frog_bram[3699] = 6'b001100;
frog_bram[3700] = 6'b001100;
frog_bram[3701] = 6'b001100;
frog_bram[3702] = 6'b110000;
frog_bram[3703] = 6'b010000;
frog_bram[3704] = 6'b010000;
frog_bram[3705] = 6'b110000;
frog_bram[3706] = 6'b001100;
frog_bram[3707] = 6'b001100;
frog_bram[3708] = 6'b001100;
frog_bram[3709] = 6'b000000;
frog_bram[3710] = 6'b000000;
frog_bram[3711] = 6'b000000;
frog_bram[3712] = 6'b000000;
frog_bram[3713] = 6'b000000;
frog_bram[3714] = 6'b000000;
frog_bram[3715] = 6'b000000;
frog_bram[3716] = 6'b000000;
frog_bram[3717] = 6'b001000;
frog_bram[3718] = 6'b001000;
frog_bram[3719] = 6'b001100;
frog_bram[3720] = 6'b001100;
frog_bram[3721] = 6'b001000;
frog_bram[3722] = 6'b001100;
frog_bram[3723] = 6'b001100;
frog_bram[3724] = 6'b001100;
frog_bram[3725] = 6'b001100;
frog_bram[3726] = 6'b001100;
frog_bram[3727] = 6'b001100;
frog_bram[3728] = 6'b001100;
frog_bram[3729] = 6'b001100;
frog_bram[3730] = 6'b001100;
frog_bram[3731] = 6'b001100;
frog_bram[3732] = 6'b001100;
frog_bram[3733] = 6'b001100;
frog_bram[3734] = 6'b110000;
frog_bram[3735] = 6'b010000;
frog_bram[3736] = 6'b010000;
frog_bram[3737] = 6'b110000;
frog_bram[3738] = 6'b001100;
frog_bram[3739] = 6'b001000;
frog_bram[3740] = 6'b000000;
frog_bram[3741] = 6'b000000;
frog_bram[3742] = 6'b000000;
frog_bram[3743] = 6'b000000;
frog_bram[3744] = 6'b000000;
frog_bram[3745] = 6'b000000;
frog_bram[3746] = 6'b000000;
frog_bram[3747] = 6'b000000;
frog_bram[3748] = 6'b000000;
frog_bram[3749] = 6'b000000;
frog_bram[3750] = 6'b000000;
frog_bram[3751] = 6'b001000;
frog_bram[3752] = 6'b001000;
frog_bram[3753] = 6'b001000;
frog_bram[3754] = 6'b001100;
frog_bram[3755] = 6'b001100;
frog_bram[3756] = 6'b001100;
frog_bram[3757] = 6'b001100;
frog_bram[3758] = 6'b001100;
frog_bram[3759] = 6'b001100;
frog_bram[3760] = 6'b001100;
frog_bram[3761] = 6'b001100;
frog_bram[3762] = 6'b001000;
frog_bram[3763] = 6'b001000;
frog_bram[3764] = 6'b001100;
frog_bram[3765] = 6'b001100;
frog_bram[3766] = 6'b001100;
frog_bram[3767] = 6'b110000;
frog_bram[3768] = 6'b110000;
frog_bram[3769] = 6'b001100;
frog_bram[3770] = 6'b001000;
frog_bram[3771] = 6'b000000;
frog_bram[3772] = 6'b000000;
frog_bram[3773] = 6'b000000;
frog_bram[3774] = 6'b000000;
frog_bram[3775] = 6'b000000;
frog_bram[3776] = 6'b000000;
frog_bram[3777] = 6'b000000;
frog_bram[3778] = 6'b000000;
frog_bram[3779] = 6'b000000;
frog_bram[3780] = 6'b001000;
frog_bram[3781] = 6'b001000;
frog_bram[3782] = 6'b001000;
frog_bram[3783] = 6'b000000;
frog_bram[3784] = 6'b000000;
frog_bram[3785] = 6'b000000;
frog_bram[3786] = 6'b001000;
frog_bram[3787] = 6'b001000;
frog_bram[3788] = 6'b001100;
frog_bram[3789] = 6'b001100;
frog_bram[3790] = 6'b001100;
frog_bram[3791] = 6'b001100;
frog_bram[3792] = 6'b001100;
frog_bram[3793] = 6'b001000;
frog_bram[3794] = 6'b000000;
frog_bram[3795] = 6'b000000;
frog_bram[3796] = 6'b001100;
frog_bram[3797] = 6'b001100;
frog_bram[3798] = 6'b001100;
frog_bram[3799] = 6'b001100;
frog_bram[3800] = 6'b001100;
frog_bram[3801] = 6'b001100;
frog_bram[3802] = 6'b000000;
frog_bram[3803] = 6'b000000;
frog_bram[3804] = 6'b000000;
frog_bram[3805] = 6'b000000;
frog_bram[3806] = 6'b000000;
frog_bram[3807] = 6'b000000;
frog_bram[3808] = 6'b000000;
frog_bram[3809] = 6'b000000;
frog_bram[3810] = 6'b001000;
frog_bram[3811] = 6'b001100;
frog_bram[3812] = 6'b001100;
frog_bram[3813] = 6'b001100;
frog_bram[3814] = 6'b001100;
frog_bram[3815] = 6'b001000;
frog_bram[3816] = 6'b001000;
frog_bram[3817] = 6'b001000;
frog_bram[3818] = 6'b000000;
frog_bram[3819] = 6'b000000;
frog_bram[3820] = 6'b000000;
frog_bram[3821] = 6'b000000;
frog_bram[3822] = 6'b001000;
frog_bram[3823] = 6'b000000;
frog_bram[3824] = 6'b000000;
frog_bram[3825] = 6'b001100;
frog_bram[3826] = 6'b001000;
frog_bram[3827] = 6'b000000;
frog_bram[3828] = 6'b000000;
frog_bram[3829] = 6'b001100;
frog_bram[3830] = 6'b001100;
frog_bram[3831] = 6'b001100;
frog_bram[3832] = 6'b001100;
frog_bram[3833] = 6'b000000;
frog_bram[3834] = 6'b000000;
frog_bram[3835] = 6'b000000;
frog_bram[3836] = 6'b000000;
frog_bram[3837] = 6'b000000;
frog_bram[3838] = 6'b000000;
frog_bram[3839] = 6'b000000;
frog_bram[3840] = 6'b000000;
frog_bram[3841] = 6'b000000;
frog_bram[3842] = 6'b001100;
frog_bram[3843] = 6'b001100;
frog_bram[3844] = 6'b001100;
frog_bram[3845] = 6'b001100;
frog_bram[3846] = 6'b001100;
frog_bram[3847] = 6'b001100;
frog_bram[3848] = 6'b001100;
frog_bram[3849] = 6'b001100;
frog_bram[3850] = 6'b001000;
frog_bram[3851] = 6'b001000;
frog_bram[3852] = 6'b001000;
frog_bram[3853] = 6'b001000;
frog_bram[3854] = 6'b000000;
frog_bram[3855] = 6'b001000;
frog_bram[3856] = 6'b001100;
frog_bram[3857] = 6'b001000;
frog_bram[3858] = 6'b001000;
frog_bram[3859] = 6'b001000;
frog_bram[3860] = 6'b000000;
frog_bram[3861] = 6'b000000;
frog_bram[3862] = 6'b000000;
frog_bram[3863] = 6'b000000;
frog_bram[3864] = 6'b000000;
frog_bram[3865] = 6'b000000;
frog_bram[3866] = 6'b000000;
frog_bram[3867] = 6'b001000;
frog_bram[3868] = 6'b001000;
frog_bram[3869] = 6'b000000;
frog_bram[3870] = 6'b000000;
frog_bram[3871] = 6'b000000;
frog_bram[3872] = 6'b000000;
frog_bram[3873] = 6'b001000;
frog_bram[3874] = 6'b001100;
frog_bram[3875] = 6'b001100;
frog_bram[3876] = 6'b001100;
frog_bram[3877] = 6'b000000;
frog_bram[3878] = 6'b001000;
frog_bram[3879] = 6'b001000;
frog_bram[3880] = 6'b001100;
frog_bram[3881] = 6'b001100;
frog_bram[3882] = 6'b001100;
frog_bram[3883] = 6'b001100;
frog_bram[3884] = 6'b001100;
frog_bram[3885] = 6'b001000;
frog_bram[3886] = 6'b000000;
frog_bram[3887] = 6'b000000;
frog_bram[3888] = 6'b001000;
frog_bram[3889] = 6'b001000;
frog_bram[3890] = 6'b001000;
frog_bram[3891] = 6'b001000;
frog_bram[3892] = 6'b000000;
frog_bram[3893] = 6'b000000;
frog_bram[3894] = 6'b000000;
frog_bram[3895] = 6'b001000;
frog_bram[3896] = 6'b000100;
frog_bram[3897] = 6'b000000;
frog_bram[3898] = 6'b001100;
frog_bram[3899] = 6'b001100;
frog_bram[3900] = 6'b001000;
frog_bram[3901] = 6'b000000;
frog_bram[3902] = 6'b000000;
frog_bram[3903] = 6'b000000;
frog_bram[3904] = 6'b000000;
frog_bram[3905] = 6'b001000;
frog_bram[3906] = 6'b001100;
frog_bram[3907] = 6'b001100;
frog_bram[3908] = 6'b001100;
frog_bram[3909] = 6'b001000;
frog_bram[3910] = 6'b000000;
frog_bram[3911] = 6'b001000;
frog_bram[3912] = 6'b001000;
frog_bram[3913] = 6'b001000;
frog_bram[3914] = 6'b001000;
frog_bram[3915] = 6'b001000;
frog_bram[3916] = 6'b001000;
frog_bram[3917] = 6'b000000;
frog_bram[3918] = 6'b000000;
frog_bram[3919] = 6'b000000;
frog_bram[3920] = 6'b000000;
frog_bram[3921] = 6'b001000;
frog_bram[3922] = 6'b001000;
frog_bram[3923] = 6'b001000;
frog_bram[3924] = 6'b001000;
frog_bram[3925] = 6'b000000;
frog_bram[3926] = 6'b001100;
frog_bram[3927] = 6'b001100;
frog_bram[3928] = 6'b000100;
frog_bram[3929] = 6'b001000;
frog_bram[3930] = 6'b001100;
frog_bram[3931] = 6'b000000;
frog_bram[3932] = 6'b000000;
frog_bram[3933] = 6'b000000;
frog_bram[3934] = 6'b000000;
frog_bram[3935] = 6'b000000;
frog_bram[3936] = 6'b000000;
frog_bram[3937] = 6'b000000;
frog_bram[3938] = 6'b001000;
frog_bram[3939] = 6'b001100;
frog_bram[3940] = 6'b001100;
frog_bram[3941] = 6'b001100;
frog_bram[3942] = 6'b001000;
frog_bram[3943] = 6'b000000;
frog_bram[3944] = 6'b000000;
frog_bram[3945] = 6'b000000;
frog_bram[3946] = 6'b000000;
frog_bram[3947] = 6'b000000;
frog_bram[3948] = 6'b000000;
frog_bram[3949] = 6'b000000;
frog_bram[3950] = 6'b000000;
frog_bram[3951] = 6'b000000;
frog_bram[3952] = 6'b000000;
frog_bram[3953] = 6'b001000;
frog_bram[3954] = 6'b001000;
frog_bram[3955] = 6'b001100;
frog_bram[3956] = 6'b001100;
frog_bram[3957] = 6'b001100;
frog_bram[3958] = 6'b001100;
frog_bram[3959] = 6'b001100;
frog_bram[3960] = 6'b001100;
frog_bram[3961] = 6'b001000;
frog_bram[3962] = 6'b000100;
frog_bram[3963] = 6'b001000;
frog_bram[3964] = 6'b001000;
frog_bram[3965] = 6'b000000;
frog_bram[3966] = 6'b000000;
frog_bram[3967] = 6'b000000;
frog_bram[3968] = 6'b000000;
frog_bram[3969] = 6'b000000;
frog_bram[3970] = 6'b001000;
frog_bram[3971] = 6'b001100;
frog_bram[3972] = 6'b001100;
frog_bram[3973] = 6'b001100;
frog_bram[3974] = 6'b001100;
frog_bram[3975] = 6'b001100;
frog_bram[3976] = 6'b001100;
frog_bram[3977] = 6'b001000;
frog_bram[3978] = 6'b000000;
frog_bram[3979] = 6'b000000;
frog_bram[3980] = 6'b000000;
frog_bram[3981] = 6'b000000;
frog_bram[3982] = 6'b000000;
frog_bram[3983] = 6'b000000;
frog_bram[3984] = 6'b000000;
frog_bram[3985] = 6'b000000;
frog_bram[3986] = 6'b001000;
frog_bram[3987] = 6'b001100;
frog_bram[3988] = 6'b001100;
frog_bram[3989] = 6'b001100;
frog_bram[3990] = 6'b001100;
frog_bram[3991] = 6'b001100;
frog_bram[3992] = 6'b001100;
frog_bram[3993] = 6'b001100;
frog_bram[3994] = 6'b001100;
frog_bram[3995] = 6'b001100;
frog_bram[3996] = 6'b001100;
frog_bram[3997] = 6'b000000;
frog_bram[3998] = 6'b000000;
frog_bram[3999] = 6'b000000;
frog_bram[4000] = 6'b000000;
frog_bram[4001] = 6'b000000;
frog_bram[4002] = 6'b001000;
frog_bram[4003] = 6'b001100;
frog_bram[4004] = 6'b001100;
frog_bram[4005] = 6'b001100;
frog_bram[4006] = 6'b001000;
frog_bram[4007] = 6'b000100;
frog_bram[4008] = 6'b001100;
frog_bram[4009] = 6'b001000;
frog_bram[4010] = 6'b000000;
frog_bram[4011] = 6'b000000;
frog_bram[4012] = 6'b000000;
frog_bram[4013] = 6'b000000;
frog_bram[4014] = 6'b000000;
frog_bram[4015] = 6'b000000;
frog_bram[4016] = 6'b000000;
frog_bram[4017] = 6'b000000;
frog_bram[4018] = 6'b000000;
frog_bram[4019] = 6'b001100;
frog_bram[4020] = 6'b001100;
frog_bram[4021] = 6'b001100;
frog_bram[4022] = 6'b001100;
frog_bram[4023] = 6'b001100;
frog_bram[4024] = 6'b001100;
frog_bram[4025] = 6'b000000;
frog_bram[4026] = 6'b000000;
frog_bram[4027] = 6'b000000;
frog_bram[4028] = 6'b000000;
frog_bram[4029] = 6'b000000;
frog_bram[4030] = 6'b000000;
frog_bram[4031] = 6'b000000;
frog_bram[4032] = 6'b000000;
frog_bram[4033] = 6'b000000;
frog_bram[4034] = 6'b000000;
frog_bram[4035] = 6'b001100;
frog_bram[4036] = 6'b001100;
frog_bram[4037] = 6'b001100;
frog_bram[4038] = 6'b001100;
frog_bram[4039] = 6'b001000;
frog_bram[4040] = 6'b000000;
frog_bram[4041] = 6'b000000;
frog_bram[4042] = 6'b000000;
frog_bram[4043] = 6'b000000;
frog_bram[4044] = 6'b000000;
frog_bram[4045] = 6'b000000;
frog_bram[4046] = 6'b000000;
frog_bram[4047] = 6'b000000;
frog_bram[4048] = 6'b000000;
frog_bram[4049] = 6'b000000;
frog_bram[4050] = 6'b000000;
frog_bram[4051] = 6'b000000;
frog_bram[4052] = 6'b000000;
frog_bram[4053] = 6'b000000;
frog_bram[4054] = 6'b000000;
frog_bram[4055] = 6'b000000;
frog_bram[4056] = 6'b000000;
frog_bram[4057] = 6'b000000;
frog_bram[4058] = 6'b000000;
frog_bram[4059] = 6'b000000;
frog_bram[4060] = 6'b000000;
frog_bram[4061] = 6'b000000;
frog_bram[4062] = 6'b000000;
frog_bram[4063] = 6'b000000;
frog_bram[4064] = 6'b000000;
frog_bram[4065] = 6'b000000;
frog_bram[4066] = 6'b000000;
frog_bram[4067] = 6'b001100;
frog_bram[4068] = 6'b001000;
frog_bram[4069] = 6'b000000;
frog_bram[4070] = 6'b001100;
frog_bram[4071] = 6'b001000;
frog_bram[4072] = 6'b000000;
frog_bram[4073] = 6'b000000;
frog_bram[4074] = 6'b000000;
frog_bram[4075] = 6'b000000;
frog_bram[4076] = 6'b000000;
frog_bram[4077] = 6'b000000;
frog_bram[4078] = 6'b000000;
frog_bram[4079] = 6'b000000;
frog_bram[4080] = 6'b000000;
frog_bram[4081] = 6'b000000;
frog_bram[4082] = 6'b000000;
frog_bram[4083] = 6'b000000;
frog_bram[4084] = 6'b000000;
frog_bram[4085] = 6'b000000;
frog_bram[4086] = 6'b000000;
frog_bram[4087] = 6'b000000;
frog_bram[4088] = 6'b000000;
frog_bram[4089] = 6'b000000;
frog_bram[4090] = 6'b000000;
frog_bram[4091] = 6'b000000;
frog_bram[4092] = 6'b000000;
frog_bram[4093] = 6'b000000;
frog_bram[4094] = 6'b000000;
frog_bram[4095] = 6'b000000;
    end

    // Calculate the base address based on the direction
    wire [11:0] base_address;  // Updated to 12 bits to handle up to 4095
    assign base_address = (direction == 2'b00) ? 12'd0 :     // Up sprite (address 0-1023)
                          (direction == 2'b01) ? 12'd1024 :  // Down sprite (address 1024-2047)
                          (direction == 2'b10) ? 12'd2048 :  // Left sprite (address 2048-3071)
                          12'd3072;                          // Right sprite (address 3072-4095)

    // Calculate the BRAM address for the current (sprite_x, sprite_y) within the selected sprite
    wire [11:0] bram_address = base_address + (sprite_y * 32) + sprite_x;

    // Output the pixel data from the BRAM based on the address
    always @(posedge clk) begin
        pixel_data <= frog_bram[bram_address];
    end

endmodule
