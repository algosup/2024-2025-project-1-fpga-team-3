module blue_car_sprite_bram (
    input wire clk,                 // Clock signal
    input wire [4:0] sprite_x,      // X coordinate within the car sprite (0-31)
    input wire [4:0] sprite_y,      // Y coordinate within the car sprite (0-31)
    output reg [5:0] pixel_data    // 6-bit pixel data
);

    // Declare a 1024x6 bit Block RAM (BRAM) for storing the 32x32 car sprite (6-bit color)
    reg [5:0] blue_car_bram [0:1023];

    // Initialize the car sprite data in BRAM
    initial begin
        blue_car_bram[0] = 6'b000000;
blue_car_bram[1] = 6'b000000;
blue_car_bram[2] = 6'b000000;
blue_car_bram[3] = 6'b000000;
blue_car_bram[4] = 6'b000000;
blue_car_bram[5] = 6'b000000;
blue_car_bram[6] = 6'b000000;
blue_car_bram[7] = 6'b000000;
blue_car_bram[8] = 6'b000000;
blue_car_bram[9] = 6'b000000;
blue_car_bram[10] = 6'b000000;
blue_car_bram[11] = 6'b000000;
blue_car_bram[12] = 6'b000000;
blue_car_bram[13] = 6'b000000;
blue_car_bram[14] = 6'b000000;
blue_car_bram[15] = 6'b000000;
blue_car_bram[16] = 6'b000000;
blue_car_bram[17] = 6'b000000;
blue_car_bram[18] = 6'b000000;
blue_car_bram[19] = 6'b000000;
blue_car_bram[20] = 6'b000000;
blue_car_bram[21] = 6'b000000;
blue_car_bram[22] = 6'b000000;
blue_car_bram[23] = 6'b000000;
blue_car_bram[24] = 6'b000000;
blue_car_bram[25] = 6'b000000;
blue_car_bram[26] = 6'b000000;
blue_car_bram[27] = 6'b000000;
blue_car_bram[28] = 6'b000000;
blue_car_bram[29] = 6'b000000;
blue_car_bram[30] = 6'b000000;
blue_car_bram[31] = 6'b000000;
blue_car_bram[32] = 6'b000000;
blue_car_bram[33] = 6'b000000;
blue_car_bram[34] = 6'b000000;
blue_car_bram[35] = 6'b000000;
blue_car_bram[36] = 6'b000000;
blue_car_bram[37] = 6'b000000;
blue_car_bram[38] = 6'b000000;
blue_car_bram[39] = 6'b000000;
blue_car_bram[40] = 6'b000000;
blue_car_bram[41] = 6'b000000;
blue_car_bram[42] = 6'b000000;
blue_car_bram[43] = 6'b000000;
blue_car_bram[44] = 6'b000000;
blue_car_bram[45] = 6'b000000;
blue_car_bram[46] = 6'b000000;
blue_car_bram[47] = 6'b000000;
blue_car_bram[48] = 6'b000000;
blue_car_bram[49] = 6'b000000;
blue_car_bram[50] = 6'b000000;
blue_car_bram[51] = 6'b000000;
blue_car_bram[52] = 6'b000000;
blue_car_bram[53] = 6'b000000;
blue_car_bram[54] = 6'b000000;
blue_car_bram[55] = 6'b000000;
blue_car_bram[56] = 6'b000000;
blue_car_bram[57] = 6'b000000;
blue_car_bram[58] = 6'b000000;
blue_car_bram[59] = 6'b000000;
blue_car_bram[60] = 6'b000000;
blue_car_bram[61] = 6'b000000;
blue_car_bram[62] = 6'b000000;
blue_car_bram[63] = 6'b000000;
blue_car_bram[64] = 6'b000000;
blue_car_bram[65] = 6'b000000;
blue_car_bram[66] = 6'b000000;
blue_car_bram[67] = 6'b000000;
blue_car_bram[68] = 6'b000000;
blue_car_bram[69] = 6'b000000;
blue_car_bram[70] = 6'b000000;
blue_car_bram[71] = 6'b000000;
blue_car_bram[72] = 6'b000000;
blue_car_bram[73] = 6'b000000;
blue_car_bram[74] = 6'b000000;
blue_car_bram[75] = 6'b000000;
blue_car_bram[76] = 6'b000000;
blue_car_bram[77] = 6'b000000;
blue_car_bram[78] = 6'b000000;
blue_car_bram[79] = 6'b000000;
blue_car_bram[80] = 6'b000000;
blue_car_bram[81] = 6'b000000;
blue_car_bram[82] = 6'b000000;
blue_car_bram[83] = 6'b000000;
blue_car_bram[84] = 6'b000000;
blue_car_bram[85] = 6'b000000;
blue_car_bram[86] = 6'b000000;
blue_car_bram[87] = 6'b000000;
blue_car_bram[88] = 6'b000000;
blue_car_bram[89] = 6'b000000;
blue_car_bram[90] = 6'b000000;
blue_car_bram[91] = 6'b000000;
blue_car_bram[92] = 6'b000000;
blue_car_bram[93] = 6'b000000;
blue_car_bram[94] = 6'b000000;
blue_car_bram[95] = 6'b000000;
blue_car_bram[96] = 6'b000000;
blue_car_bram[97] = 6'b000000;
blue_car_bram[98] = 6'b000000;
blue_car_bram[99] = 6'b000000;
blue_car_bram[100] = 6'b000000;
blue_car_bram[101] = 6'b000000;
blue_car_bram[102] = 6'b000000;
blue_car_bram[103] = 6'b000000;
blue_car_bram[104] = 6'b000000;
blue_car_bram[105] = 6'b000000;
blue_car_bram[106] = 6'b000000;
blue_car_bram[107] = 6'b000000;
blue_car_bram[108] = 6'b000000;
blue_car_bram[109] = 6'b000000;
blue_car_bram[110] = 6'b000000;
blue_car_bram[111] = 6'b000000;
blue_car_bram[112] = 6'b000000;
blue_car_bram[113] = 6'b000000;
blue_car_bram[114] = 6'b000000;
blue_car_bram[115] = 6'b000000;
blue_car_bram[116] = 6'b000000;
blue_car_bram[117] = 6'b000000;
blue_car_bram[118] = 6'b000000;
blue_car_bram[119] = 6'b000000;
blue_car_bram[120] = 6'b000000;
blue_car_bram[121] = 6'b000000;
blue_car_bram[122] = 6'b000000;
blue_car_bram[123] = 6'b000000;
blue_car_bram[124] = 6'b000000;
blue_car_bram[125] = 6'b000000;
blue_car_bram[126] = 6'b000000;
blue_car_bram[127] = 6'b000000;
blue_car_bram[128] = 6'b000000;
blue_car_bram[129] = 6'b000000;
blue_car_bram[130] = 6'b000000;
blue_car_bram[131] = 6'b000000;
blue_car_bram[132] = 6'b000000;
blue_car_bram[133] = 6'b000000;
blue_car_bram[134] = 6'b010101;
blue_car_bram[135] = 6'b010101;
blue_car_bram[136] = 6'b010101;
blue_car_bram[137] = 6'b010101;
blue_car_bram[138] = 6'b010101;
blue_car_bram[139] = 6'b010101;
blue_car_bram[140] = 6'b000000;
blue_car_bram[141] = 6'b000000;
blue_car_bram[142] = 6'b000000;
blue_car_bram[143] = 6'b000000;
blue_car_bram[144] = 6'b000000;
blue_car_bram[145] = 6'b000000;
blue_car_bram[146] = 6'b000000;
blue_car_bram[147] = 6'b000000;
blue_car_bram[148] = 6'b010101;
blue_car_bram[149] = 6'b010101;
blue_car_bram[150] = 6'b010101;
blue_car_bram[151] = 6'b010101;
blue_car_bram[152] = 6'b010101;
blue_car_bram[153] = 6'b010101;
blue_car_bram[154] = 6'b000000;
blue_car_bram[155] = 6'b000000;
blue_car_bram[156] = 6'b000000;
blue_car_bram[157] = 6'b000000;
blue_car_bram[158] = 6'b000000;
blue_car_bram[159] = 6'b000000;
blue_car_bram[160] = 6'b000000;
blue_car_bram[161] = 6'b000000;
blue_car_bram[162] = 6'b000000;
blue_car_bram[163] = 6'b000000;
blue_car_bram[164] = 6'b000000;
blue_car_bram[165] = 6'b010101;
blue_car_bram[166] = 6'b010101;
blue_car_bram[167] = 6'b010101;
blue_car_bram[168] = 6'b010101;
blue_car_bram[169] = 6'b010101;
blue_car_bram[170] = 6'b010101;
blue_car_bram[171] = 6'b010101;
blue_car_bram[172] = 6'b010101;
blue_car_bram[173] = 6'b000000;
blue_car_bram[174] = 6'b000000;
blue_car_bram[175] = 6'b000000;
blue_car_bram[176] = 6'b000000;
blue_car_bram[177] = 6'b000000;
blue_car_bram[178] = 6'b000000;
blue_car_bram[179] = 6'b010101;
blue_car_bram[180] = 6'b010101;
blue_car_bram[181] = 6'b010101;
blue_car_bram[182] = 6'b010101;
blue_car_bram[183] = 6'b010101;
blue_car_bram[184] = 6'b010101;
blue_car_bram[185] = 6'b010101;
blue_car_bram[186] = 6'b010101;
blue_car_bram[187] = 6'b000000;
blue_car_bram[188] = 6'b000000;
blue_car_bram[189] = 6'b000000;
blue_car_bram[190] = 6'b000000;
blue_car_bram[191] = 6'b000000;
blue_car_bram[192] = 6'b000000;
blue_car_bram[193] = 6'b000000;
blue_car_bram[194] = 6'b000000;
blue_car_bram[195] = 6'b000000;
blue_car_bram[196] = 6'b000000;
blue_car_bram[197] = 6'b000000;
blue_car_bram[198] = 6'b000000;
blue_car_bram[199] = 6'b000000;
blue_car_bram[200] = 6'b000000;
blue_car_bram[201] = 6'b000000;
blue_car_bram[202] = 6'b000000;
blue_car_bram[203] = 6'b000000;
blue_car_bram[204] = 6'b000000;
blue_car_bram[205] = 6'b000000;
blue_car_bram[206] = 6'b000000;
blue_car_bram[207] = 6'b000000;
blue_car_bram[208] = 6'b000000;
blue_car_bram[209] = 6'b000000;
blue_car_bram[210] = 6'b000000;
blue_car_bram[211] = 6'b000000;
blue_car_bram[212] = 6'b000000;
blue_car_bram[213] = 6'b000000;
blue_car_bram[214] = 6'b000000;
blue_car_bram[215] = 6'b000000;
blue_car_bram[216] = 6'b000000;
blue_car_bram[217] = 6'b000000;
blue_car_bram[218] = 6'b000000;
blue_car_bram[219] = 6'b000000;
blue_car_bram[220] = 6'b000000;
blue_car_bram[221] = 6'b000000;
blue_car_bram[222] = 6'b000000;
blue_car_bram[223] = 6'b000000;
blue_car_bram[224] = 6'b000000;
blue_car_bram[225] = 6'b000000;
blue_car_bram[226] = 6'b101001;
blue_car_bram[227] = 6'b000000;
blue_car_bram[228] = 6'b000110;
blue_car_bram[229] = 6'b000110;
blue_car_bram[230] = 6'b000110;
blue_car_bram[231] = 6'b000110;
blue_car_bram[232] = 6'b000110;
blue_car_bram[233] = 6'b000110;
blue_car_bram[234] = 6'b000110;
blue_car_bram[235] = 6'b000110;
blue_car_bram[236] = 6'b000110;
blue_car_bram[237] = 6'b000110;
blue_car_bram[238] = 6'b000110;
blue_car_bram[239] = 6'b000110;
blue_car_bram[240] = 6'b000110;
blue_car_bram[241] = 6'b000110;
blue_car_bram[242] = 6'b000110;
blue_car_bram[243] = 6'b000110;
blue_car_bram[244] = 6'b000110;
blue_car_bram[245] = 6'b000110;
blue_car_bram[246] = 6'b000110;
blue_car_bram[247] = 6'b000110;
blue_car_bram[248] = 6'b000110;
blue_car_bram[249] = 6'b000110;
blue_car_bram[250] = 6'b000110;
blue_car_bram[251] = 6'b000110;
blue_car_bram[252] = 6'b000110;
blue_car_bram[253] = 6'b000000;
blue_car_bram[254] = 6'b000000;
blue_car_bram[255] = 6'b000000;
blue_car_bram[256] = 6'b000000;
blue_car_bram[257] = 6'b101001;
blue_car_bram[258] = 6'b111101;
blue_car_bram[259] = 6'b000000;
blue_car_bram[260] = 6'b000111;
blue_car_bram[261] = 6'b000111;
blue_car_bram[262] = 6'b000000;
blue_car_bram[263] = 6'b000000;
blue_car_bram[264] = 6'b000000;
blue_car_bram[265] = 6'b000000;
blue_car_bram[266] = 6'b000000;
blue_car_bram[267] = 6'b000000;
blue_car_bram[268] = 6'b000000;
blue_car_bram[269] = 6'b000000;
blue_car_bram[270] = 6'b000000;
blue_car_bram[271] = 6'b000111;
blue_car_bram[272] = 6'b000111;
blue_car_bram[273] = 6'b000000;
blue_car_bram[274] = 6'b000000;
blue_car_bram[275] = 6'b000000;
blue_car_bram[276] = 6'b000000;
blue_car_bram[277] = 6'b000000;
blue_car_bram[278] = 6'b000000;
blue_car_bram[279] = 6'b000000;
blue_car_bram[280] = 6'b000000;
blue_car_bram[281] = 6'b000000;
blue_car_bram[282] = 6'b000000;
blue_car_bram[283] = 6'b000111;
blue_car_bram[284] = 6'b000111;
blue_car_bram[285] = 6'b000010;
blue_car_bram[286] = 6'b000000;
blue_car_bram[287] = 6'b000000;
blue_car_bram[288] = 6'b000000;
blue_car_bram[289] = 6'b101001;
blue_car_bram[290] = 6'b000000;
blue_car_bram[291] = 6'b000010;
blue_car_bram[292] = 6'b000011;
blue_car_bram[293] = 6'b000111;
blue_car_bram[294] = 6'b000110;
blue_car_bram[295] = 6'b000110;
blue_car_bram[296] = 6'b000000;
blue_car_bram[297] = 6'b000000;
blue_car_bram[298] = 6'b000000;
blue_car_bram[299] = 6'b000000;
blue_car_bram[300] = 6'b000000;
blue_car_bram[301] = 6'b000000;
blue_car_bram[302] = 6'b000000;
blue_car_bram[303] = 6'b000111;
blue_car_bram[304] = 6'b000111;
blue_car_bram[305] = 6'b000000;
blue_car_bram[306] = 6'b000000;
blue_car_bram[307] = 6'b000000;
blue_car_bram[308] = 6'b000000;
blue_car_bram[309] = 6'b000000;
blue_car_bram[310] = 6'b000000;
blue_car_bram[311] = 6'b000000;
blue_car_bram[312] = 6'b000000;
blue_car_bram[313] = 6'b000110;
blue_car_bram[314] = 6'b000110;
blue_car_bram[315] = 6'b000111;
blue_car_bram[316] = 6'b000111;
blue_car_bram[317] = 6'b000011;
blue_car_bram[318] = 6'b000000;
blue_car_bram[319] = 6'b000000;
blue_car_bram[320] = 6'b000000;
blue_car_bram[321] = 6'b000000;
blue_car_bram[322] = 6'b000010;
blue_car_bram[323] = 6'b000011;
blue_car_bram[324] = 6'b000000;
blue_car_bram[325] = 6'b000000;
blue_car_bram[326] = 6'b000111;
blue_car_bram[327] = 6'b000111;
blue_car_bram[328] = 6'b000110;
blue_car_bram[329] = 6'b000110;
blue_car_bram[330] = 6'b000110;
blue_car_bram[331] = 6'b000110;
blue_car_bram[332] = 6'b000110;
blue_car_bram[333] = 6'b000110;
blue_car_bram[334] = 6'b000110;
blue_car_bram[335] = 6'b000111;
blue_car_bram[336] = 6'b000111;
blue_car_bram[337] = 6'b000110;
blue_car_bram[338] = 6'b000110;
blue_car_bram[339] = 6'b000110;
blue_car_bram[340] = 6'b000110;
blue_car_bram[341] = 6'b000110;
blue_car_bram[342] = 6'b000110;
blue_car_bram[343] = 6'b000110;
blue_car_bram[344] = 6'b000110;
blue_car_bram[345] = 6'b000111;
blue_car_bram[346] = 6'b000111;
blue_car_bram[347] = 6'b000111;
blue_car_bram[348] = 6'b000011;
blue_car_bram[349] = 6'b000000;
blue_car_bram[350] = 6'b100101;
blue_car_bram[351] = 6'b000000;
blue_car_bram[352] = 6'b000000;
blue_car_bram[353] = 6'b000000;
blue_car_bram[354] = 6'b000011;
blue_car_bram[355] = 6'b000000;
blue_car_bram[356] = 6'b000000;
blue_car_bram[357] = 6'b000000;
blue_car_bram[358] = 6'b000000;
blue_car_bram[359] = 6'b000000;
blue_car_bram[360] = 6'b000111;
blue_car_bram[361] = 6'b000111;
blue_car_bram[362] = 6'b000111;
blue_car_bram[363] = 6'b000001;
blue_car_bram[364] = 6'b000111;
blue_car_bram[365] = 6'b000111;
blue_car_bram[366] = 6'b000111;
blue_car_bram[367] = 6'b000111;
blue_car_bram[368] = 6'b000111;
blue_car_bram[369] = 6'b000111;
blue_car_bram[370] = 6'b000111;
blue_car_bram[371] = 6'b000111;
blue_car_bram[372] = 6'b000111;
blue_car_bram[373] = 6'b000111;
blue_car_bram[374] = 6'b000001;
blue_car_bram[375] = 6'b000111;
blue_car_bram[376] = 6'b000111;
blue_car_bram[377] = 6'b000011;
blue_car_bram[378] = 6'b000000;
blue_car_bram[379] = 6'b000000;
blue_car_bram[380] = 6'b000010;
blue_car_bram[381] = 6'b000000;
blue_car_bram[382] = 6'b100101;
blue_car_bram[383] = 6'b000000;
blue_car_bram[384] = 6'b000000;
blue_car_bram[385] = 6'b000001;
blue_car_bram[386] = 6'b000011;
blue_car_bram[387] = 6'b000000;
blue_car_bram[388] = 6'b000000;
blue_car_bram[389] = 6'b000000;
blue_car_bram[390] = 6'b101010;
blue_car_bram[391] = 6'b000000;
blue_car_bram[392] = 6'b000000;
blue_car_bram[393] = 6'b000011;
blue_car_bram[394] = 6'b000001;
blue_car_bram[395] = 6'b000010;
blue_car_bram[396] = 6'b000011;
blue_car_bram[397] = 6'b000011;
blue_car_bram[398] = 6'b000011;
blue_car_bram[399] = 6'b000111;
blue_car_bram[400] = 6'b000111;
blue_car_bram[401] = 6'b000011;
blue_car_bram[402] = 6'b000011;
blue_car_bram[403] = 6'b000011;
blue_car_bram[404] = 6'b000011;
blue_car_bram[405] = 6'b000011;
blue_car_bram[406] = 6'b000010;
blue_car_bram[407] = 6'b000001;
blue_car_bram[408] = 6'b000011;
blue_car_bram[409] = 6'b000000;
blue_car_bram[410] = 6'b000000;
blue_car_bram[411] = 6'b000000;
blue_car_bram[412] = 6'b000011;
blue_car_bram[413] = 6'b000010;
blue_car_bram[414] = 6'b000000;
blue_car_bram[415] = 6'b000000;
blue_car_bram[416] = 6'b000000;
blue_car_bram[417] = 6'b000001;
blue_car_bram[418] = 6'b000011;
blue_car_bram[419] = 6'b000000;
blue_car_bram[420] = 6'b000000;
blue_car_bram[421] = 6'b101010;
blue_car_bram[422] = 6'b000000;
blue_car_bram[423] = 6'b000000;
blue_car_bram[424] = 6'b000000;
blue_car_bram[425] = 6'b000011;
blue_car_bram[426] = 6'b000010;
blue_car_bram[427] = 6'b000111;
blue_car_bram[428] = 6'b000111;
blue_car_bram[429] = 6'b000111;
blue_car_bram[430] = 6'b000111;
blue_car_bram[431] = 6'b000111;
blue_car_bram[432] = 6'b000111;
blue_car_bram[433] = 6'b000111;
blue_car_bram[434] = 6'b000111;
blue_car_bram[435] = 6'b000111;
blue_car_bram[436] = 6'b000111;
blue_car_bram[437] = 6'b000111;
blue_car_bram[438] = 6'b000111;
blue_car_bram[439] = 6'b000010;
blue_car_bram[440] = 6'b000011;
blue_car_bram[441] = 6'b000000;
blue_car_bram[442] = 6'b000000;
blue_car_bram[443] = 6'b000000;
blue_car_bram[444] = 6'b000111;
blue_car_bram[445] = 6'b101111;
blue_car_bram[446] = 6'b000000;
blue_car_bram[447] = 6'b000000;
blue_car_bram[448] = 6'b000000;
blue_car_bram[449] = 6'b000001;
blue_car_bram[450] = 6'b000011;
blue_car_bram[451] = 6'b000000;
blue_car_bram[452] = 6'b000000;
blue_car_bram[453] = 6'b000000;
blue_car_bram[454] = 6'b000000;
blue_car_bram[455] = 6'b000000;
blue_car_bram[456] = 6'b000000;
blue_car_bram[457] = 6'b000011;
blue_car_bram[458] = 6'b000111;
blue_car_bram[459] = 6'b000111;
blue_car_bram[460] = 6'b000111;
blue_car_bram[461] = 6'b000111;
blue_car_bram[462] = 6'b000111;
blue_car_bram[463] = 6'b000111;
blue_car_bram[464] = 6'b000111;
blue_car_bram[465] = 6'b000111;
blue_car_bram[466] = 6'b000111;
blue_car_bram[467] = 6'b000111;
blue_car_bram[468] = 6'b000111;
blue_car_bram[469] = 6'b000111;
blue_car_bram[470] = 6'b000111;
blue_car_bram[471] = 6'b000111;
blue_car_bram[472] = 6'b000011;
blue_car_bram[473] = 6'b000000;
blue_car_bram[474] = 6'b000000;
blue_car_bram[475] = 6'b000000;
blue_car_bram[476] = 6'b000111;
blue_car_bram[477] = 6'b111111;
blue_car_bram[478] = 6'b000000;
blue_car_bram[479] = 6'b000000;
blue_car_bram[480] = 6'b000000;
blue_car_bram[481] = 6'b000001;
blue_car_bram[482] = 6'b000011;
blue_car_bram[483] = 6'b000000;
blue_car_bram[484] = 6'b000000;
blue_car_bram[485] = 6'b000000;
blue_car_bram[486] = 6'b000000;
blue_car_bram[487] = 6'b000000;
blue_car_bram[488] = 6'b000000;
blue_car_bram[489] = 6'b000011;
blue_car_bram[490] = 6'b000111;
blue_car_bram[491] = 6'b000111;
blue_car_bram[492] = 6'b000111;
blue_car_bram[493] = 6'b000111;
blue_car_bram[494] = 6'b000111;
blue_car_bram[495] = 6'b000111;
blue_car_bram[496] = 6'b000111;
blue_car_bram[497] = 6'b000111;
blue_car_bram[498] = 6'b000111;
blue_car_bram[499] = 6'b000111;
blue_car_bram[500] = 6'b000111;
blue_car_bram[501] = 6'b000111;
blue_car_bram[502] = 6'b000111;
blue_car_bram[503] = 6'b000111;
blue_car_bram[504] = 6'b000011;
blue_car_bram[505] = 6'b000000;
blue_car_bram[506] = 6'b000000;
blue_car_bram[507] = 6'b000000;
blue_car_bram[508] = 6'b000111;
blue_car_bram[509] = 6'b111111;
blue_car_bram[510] = 6'b000000;
blue_car_bram[511] = 6'b000000;
blue_car_bram[512] = 6'b000000;
blue_car_bram[513] = 6'b000001;
blue_car_bram[514] = 6'b000011;
blue_car_bram[515] = 6'b000000;
blue_car_bram[516] = 6'b000000;
blue_car_bram[517] = 6'b000000;
blue_car_bram[518] = 6'b000000;
blue_car_bram[519] = 6'b000000;
blue_car_bram[520] = 6'b000000;
blue_car_bram[521] = 6'b000011;
blue_car_bram[522] = 6'b000111;
blue_car_bram[523] = 6'b000111;
blue_car_bram[524] = 6'b000111;
blue_car_bram[525] = 6'b000111;
blue_car_bram[526] = 6'b000111;
blue_car_bram[527] = 6'b000111;
blue_car_bram[528] = 6'b000111;
blue_car_bram[529] = 6'b000111;
blue_car_bram[530] = 6'b000111;
blue_car_bram[531] = 6'b000111;
blue_car_bram[532] = 6'b000111;
blue_car_bram[533] = 6'b000111;
blue_car_bram[534] = 6'b000111;
blue_car_bram[535] = 6'b000111;
blue_car_bram[536] = 6'b000011;
blue_car_bram[537] = 6'b000000;
blue_car_bram[538] = 6'b000000;
blue_car_bram[539] = 6'b000000;
blue_car_bram[540] = 6'b000111;
blue_car_bram[541] = 6'b111111;
blue_car_bram[542] = 6'b000000;
blue_car_bram[543] = 6'b000000;
blue_car_bram[544] = 6'b000000;
blue_car_bram[545] = 6'b000001;
blue_car_bram[546] = 6'b000011;
blue_car_bram[547] = 6'b000000;
blue_car_bram[548] = 6'b000000;
blue_car_bram[549] = 6'b000000;
blue_car_bram[550] = 6'b101010;
blue_car_bram[551] = 6'b000000;
blue_car_bram[552] = 6'b000000;
blue_car_bram[553] = 6'b000011;
blue_car_bram[554] = 6'b000111;
blue_car_bram[555] = 6'b000111;
blue_car_bram[556] = 6'b000111;
blue_car_bram[557] = 6'b000111;
blue_car_bram[558] = 6'b000111;
blue_car_bram[559] = 6'b000111;
blue_car_bram[560] = 6'b000111;
blue_car_bram[561] = 6'b000111;
blue_car_bram[562] = 6'b000111;
blue_car_bram[563] = 6'b000111;
blue_car_bram[564] = 6'b000111;
blue_car_bram[565] = 6'b000111;
blue_car_bram[566] = 6'b000111;
blue_car_bram[567] = 6'b000111;
blue_car_bram[568] = 6'b000011;
blue_car_bram[569] = 6'b000000;
blue_car_bram[570] = 6'b000000;
blue_car_bram[571] = 6'b000000;
blue_car_bram[572] = 6'b000111;
blue_car_bram[573] = 6'b111111;
blue_car_bram[574] = 6'b000000;
blue_car_bram[575] = 6'b000000;
blue_car_bram[576] = 6'b000000;
blue_car_bram[577] = 6'b000001;
blue_car_bram[578] = 6'b000011;
blue_car_bram[579] = 6'b000000;
blue_car_bram[580] = 6'b000000;
blue_car_bram[581] = 6'b101010;
blue_car_bram[582] = 6'b000000;
blue_car_bram[583] = 6'b000000;
blue_car_bram[584] = 6'b000000;
blue_car_bram[585] = 6'b000010;
blue_car_bram[586] = 6'b000001;
blue_car_bram[587] = 6'b000011;
blue_car_bram[588] = 6'b000111;
blue_car_bram[589] = 6'b000111;
blue_car_bram[590] = 6'b000111;
blue_car_bram[591] = 6'b000111;
blue_car_bram[592] = 6'b000111;
blue_car_bram[593] = 6'b000111;
blue_car_bram[594] = 6'b000111;
blue_car_bram[595] = 6'b000111;
blue_car_bram[596] = 6'b000111;
blue_car_bram[597] = 6'b000111;
blue_car_bram[598] = 6'b000011;
blue_car_bram[599] = 6'b000001;
blue_car_bram[600] = 6'b000010;
blue_car_bram[601] = 6'b000000;
blue_car_bram[602] = 6'b000000;
blue_car_bram[603] = 6'b000000;
blue_car_bram[604] = 6'b000011;
blue_car_bram[605] = 6'b000111;
blue_car_bram[606] = 6'b000000;
blue_car_bram[607] = 6'b000000;
blue_car_bram[608] = 6'b000000;
blue_car_bram[609] = 6'b000001;
blue_car_bram[610] = 6'b000011;
blue_car_bram[611] = 6'b000000;
blue_car_bram[612] = 6'b000000;
blue_car_bram[613] = 6'b000000;
blue_car_bram[614] = 6'b000000;
blue_car_bram[615] = 6'b000000;
blue_car_bram[616] = 6'b000010;
blue_car_bram[617] = 6'b000111;
blue_car_bram[618] = 6'b000010;
blue_car_bram[619] = 6'b000001;
blue_car_bram[620] = 6'b000011;
blue_car_bram[621] = 6'b000111;
blue_car_bram[622] = 6'b000111;
blue_car_bram[623] = 6'b000111;
blue_car_bram[624] = 6'b000111;
blue_car_bram[625] = 6'b000111;
blue_car_bram[626] = 6'b000111;
blue_car_bram[627] = 6'b000111;
blue_car_bram[628] = 6'b000111;
blue_car_bram[629] = 6'b000011;
blue_car_bram[630] = 6'b000001;
blue_car_bram[631] = 6'b000010;
blue_car_bram[632] = 6'b000111;
blue_car_bram[633] = 6'b000010;
blue_car_bram[634] = 6'b000000;
blue_car_bram[635] = 6'b000000;
blue_car_bram[636] = 6'b000010;
blue_car_bram[637] = 6'b000000;
blue_car_bram[638] = 6'b100101;
blue_car_bram[639] = 6'b000000;
blue_car_bram[640] = 6'b000000;
blue_car_bram[641] = 6'b000000;
blue_car_bram[642] = 6'b000011;
blue_car_bram[643] = 6'b000010;
blue_car_bram[644] = 6'b000000;
blue_car_bram[645] = 6'b000000;
blue_car_bram[646] = 6'b000010;
blue_car_bram[647] = 6'b000010;
blue_car_bram[648] = 6'b000111;
blue_car_bram[649] = 6'b000111;
blue_car_bram[650] = 6'b000111;
blue_car_bram[651] = 6'b000110;
blue_car_bram[652] = 6'b000111;
blue_car_bram[653] = 6'b000111;
blue_car_bram[654] = 6'b000111;
blue_car_bram[655] = 6'b000111;
blue_car_bram[656] = 6'b000111;
blue_car_bram[657] = 6'b000111;
blue_car_bram[658] = 6'b000111;
blue_car_bram[659] = 6'b000111;
blue_car_bram[660] = 6'b000111;
blue_car_bram[661] = 6'b000111;
blue_car_bram[662] = 6'b000110;
blue_car_bram[663] = 6'b000111;
blue_car_bram[664] = 6'b000111;
blue_car_bram[665] = 6'b000111;
blue_car_bram[666] = 6'b000010;
blue_car_bram[667] = 6'b000010;
blue_car_bram[668] = 6'b000011;
blue_car_bram[669] = 6'b000000;
blue_car_bram[670] = 6'b100101;
blue_car_bram[671] = 6'b000000;
blue_car_bram[672] = 6'b000000;
blue_car_bram[673] = 6'b101001;
blue_car_bram[674] = 6'b000001;
blue_car_bram[675] = 6'b000011;
blue_car_bram[676] = 6'b000010;
blue_car_bram[677] = 6'b000010;
blue_car_bram[678] = 6'b000111;
blue_car_bram[679] = 6'b000111;
blue_car_bram[680] = 6'b000000;
blue_car_bram[681] = 6'b000000;
blue_car_bram[682] = 6'b000000;
blue_car_bram[683] = 6'b000000;
blue_car_bram[684] = 6'b000000;
blue_car_bram[685] = 6'b000000;
blue_car_bram[686] = 6'b000000;
blue_car_bram[687] = 6'b000111;
blue_car_bram[688] = 6'b000111;
blue_car_bram[689] = 6'b000000;
blue_car_bram[690] = 6'b000000;
blue_car_bram[691] = 6'b000000;
blue_car_bram[692] = 6'b000000;
blue_car_bram[693] = 6'b000000;
blue_car_bram[694] = 6'b000000;
blue_car_bram[695] = 6'b000000;
blue_car_bram[696] = 6'b000000;
blue_car_bram[697] = 6'b000111;
blue_car_bram[698] = 6'b000111;
blue_car_bram[699] = 6'b000111;
blue_car_bram[700] = 6'b000011;
blue_car_bram[701] = 6'b000010;
blue_car_bram[702] = 6'b000000;
blue_car_bram[703] = 6'b000000;
blue_car_bram[704] = 6'b000000;
blue_car_bram[705] = 6'b111101;
blue_car_bram[706] = 6'b101001;
blue_car_bram[707] = 6'b000000;
blue_car_bram[708] = 6'b000011;
blue_car_bram[709] = 6'b000111;
blue_car_bram[710] = 6'b000000;
blue_car_bram[711] = 6'b000000;
blue_car_bram[712] = 6'b000000;
blue_car_bram[713] = 6'b000000;
blue_car_bram[714] = 6'b000000;
blue_car_bram[715] = 6'b000000;
blue_car_bram[716] = 6'b000000;
blue_car_bram[717] = 6'b000000;
blue_car_bram[718] = 6'b000000;
blue_car_bram[719] = 6'b000111;
blue_car_bram[720] = 6'b000111;
blue_car_bram[721] = 6'b000000;
blue_car_bram[722] = 6'b000000;
blue_car_bram[723] = 6'b000000;
blue_car_bram[724] = 6'b000000;
blue_car_bram[725] = 6'b000000;
blue_car_bram[726] = 6'b000000;
blue_car_bram[727] = 6'b000000;
blue_car_bram[728] = 6'b000000;
blue_car_bram[729] = 6'b000000;
blue_car_bram[730] = 6'b000000;
blue_car_bram[731] = 6'b000111;
blue_car_bram[732] = 6'b000111;
blue_car_bram[733] = 6'b000011;
blue_car_bram[734] = 6'b000000;
blue_car_bram[735] = 6'b000000;
blue_car_bram[736] = 6'b000000;
blue_car_bram[737] = 6'b000000;
blue_car_bram[738] = 6'b111101;
blue_car_bram[739] = 6'b000000;
blue_car_bram[740] = 6'b000111;
blue_car_bram[741] = 6'b000111;
blue_car_bram[742] = 6'b000110;
blue_car_bram[743] = 6'b000110;
blue_car_bram[744] = 6'b000110;
blue_car_bram[745] = 6'b000110;
blue_car_bram[746] = 6'b000110;
blue_car_bram[747] = 6'b000110;
blue_car_bram[748] = 6'b000110;
blue_car_bram[749] = 6'b000110;
blue_car_bram[750] = 6'b000110;
blue_car_bram[751] = 6'b000111;
blue_car_bram[752] = 6'b000111;
blue_car_bram[753] = 6'b000110;
blue_car_bram[754] = 6'b000110;
blue_car_bram[755] = 6'b000110;
blue_car_bram[756] = 6'b000110;
blue_car_bram[757] = 6'b000110;
blue_car_bram[758] = 6'b000110;
blue_car_bram[759] = 6'b000110;
blue_car_bram[760] = 6'b000110;
blue_car_bram[761] = 6'b000110;
blue_car_bram[762] = 6'b000110;
blue_car_bram[763] = 6'b000111;
blue_car_bram[764] = 6'b000111;
blue_car_bram[765] = 6'b000000;
blue_car_bram[766] = 6'b000000;
blue_car_bram[767] = 6'b000000;
blue_car_bram[768] = 6'b000000;
blue_car_bram[769] = 6'b000000;
blue_car_bram[770] = 6'b000000;
blue_car_bram[771] = 6'b000000;
blue_car_bram[772] = 6'b000000;
blue_car_bram[773] = 6'b000000;
blue_car_bram[774] = 6'b000000;
blue_car_bram[775] = 6'b000000;
blue_car_bram[776] = 6'b000000;
blue_car_bram[777] = 6'b000000;
blue_car_bram[778] = 6'b000000;
blue_car_bram[779] = 6'b000000;
blue_car_bram[780] = 6'b000000;
blue_car_bram[781] = 6'b000000;
blue_car_bram[782] = 6'b000000;
blue_car_bram[783] = 6'b000000;
blue_car_bram[784] = 6'b000000;
blue_car_bram[785] = 6'b000000;
blue_car_bram[786] = 6'b000000;
blue_car_bram[787] = 6'b000000;
blue_car_bram[788] = 6'b000000;
blue_car_bram[789] = 6'b000000;
blue_car_bram[790] = 6'b000000;
blue_car_bram[791] = 6'b000000;
blue_car_bram[792] = 6'b000000;
blue_car_bram[793] = 6'b000000;
blue_car_bram[794] = 6'b000000;
blue_car_bram[795] = 6'b000000;
blue_car_bram[796] = 6'b000000;
blue_car_bram[797] = 6'b000000;
blue_car_bram[798] = 6'b000000;
blue_car_bram[799] = 6'b000000;
blue_car_bram[800] = 6'b000000;
blue_car_bram[801] = 6'b000000;
blue_car_bram[802] = 6'b000000;
blue_car_bram[803] = 6'b000000;
blue_car_bram[804] = 6'b000000;
blue_car_bram[805] = 6'b010101;
blue_car_bram[806] = 6'b000000;
blue_car_bram[807] = 6'b000000;
blue_car_bram[808] = 6'b000000;
blue_car_bram[809] = 6'b000000;
blue_car_bram[810] = 6'b000000;
blue_car_bram[811] = 6'b000000;
blue_car_bram[812] = 6'b010101;
blue_car_bram[813] = 6'b000000;
blue_car_bram[814] = 6'b000000;
blue_car_bram[815] = 6'b000000;
blue_car_bram[816] = 6'b000000;
blue_car_bram[817] = 6'b000000;
blue_car_bram[818] = 6'b000000;
blue_car_bram[819] = 6'b010101;
blue_car_bram[820] = 6'b000000;
blue_car_bram[821] = 6'b000000;
blue_car_bram[822] = 6'b000000;
blue_car_bram[823] = 6'b000000;
blue_car_bram[824] = 6'b000000;
blue_car_bram[825] = 6'b000000;
blue_car_bram[826] = 6'b010101;
blue_car_bram[827] = 6'b000000;
blue_car_bram[828] = 6'b000000;
blue_car_bram[829] = 6'b000000;
blue_car_bram[830] = 6'b000000;
blue_car_bram[831] = 6'b000000;
blue_car_bram[832] = 6'b000000;
blue_car_bram[833] = 6'b000000;
blue_car_bram[834] = 6'b000000;
blue_car_bram[835] = 6'b000000;
blue_car_bram[836] = 6'b000000;
blue_car_bram[837] = 6'b000000;
blue_car_bram[838] = 6'b010101;
blue_car_bram[839] = 6'b010101;
blue_car_bram[840] = 6'b010101;
blue_car_bram[841] = 6'b010101;
blue_car_bram[842] = 6'b010101;
blue_car_bram[843] = 6'b010101;
blue_car_bram[844] = 6'b000000;
blue_car_bram[845] = 6'b000000;
blue_car_bram[846] = 6'b000000;
blue_car_bram[847] = 6'b000000;
blue_car_bram[848] = 6'b000000;
blue_car_bram[849] = 6'b000000;
blue_car_bram[850] = 6'b000000;
blue_car_bram[851] = 6'b000000;
blue_car_bram[852] = 6'b010101;
blue_car_bram[853] = 6'b010101;
blue_car_bram[854] = 6'b010101;
blue_car_bram[855] = 6'b010101;
blue_car_bram[856] = 6'b010101;
blue_car_bram[857] = 6'b010101;
blue_car_bram[858] = 6'b000000;
blue_car_bram[859] = 6'b000000;
blue_car_bram[860] = 6'b000000;
blue_car_bram[861] = 6'b000000;
blue_car_bram[862] = 6'b000000;
blue_car_bram[863] = 6'b000000;
blue_car_bram[864] = 6'b000000;
blue_car_bram[865] = 6'b000000;
blue_car_bram[866] = 6'b000000;
blue_car_bram[867] = 6'b000000;
blue_car_bram[868] = 6'b000000;
blue_car_bram[869] = 6'b000000;
blue_car_bram[870] = 6'b000000;
blue_car_bram[871] = 6'b000000;
blue_car_bram[872] = 6'b000000;
blue_car_bram[873] = 6'b000000;
blue_car_bram[874] = 6'b000000;
blue_car_bram[875] = 6'b000000;
blue_car_bram[876] = 6'b000000;
blue_car_bram[877] = 6'b000000;
blue_car_bram[878] = 6'b000000;
blue_car_bram[879] = 6'b000000;
blue_car_bram[880] = 6'b000000;
blue_car_bram[881] = 6'b000000;
blue_car_bram[882] = 6'b000000;
blue_car_bram[883] = 6'b000000;
blue_car_bram[884] = 6'b000000;
blue_car_bram[885] = 6'b000000;
blue_car_bram[886] = 6'b000000;
blue_car_bram[887] = 6'b000000;
blue_car_bram[888] = 6'b000000;
blue_car_bram[889] = 6'b000000;
blue_car_bram[890] = 6'b000000;
blue_car_bram[891] = 6'b000000;
blue_car_bram[892] = 6'b000000;
blue_car_bram[893] = 6'b000000;
blue_car_bram[894] = 6'b000000;
blue_car_bram[895] = 6'b000000;
blue_car_bram[896] = 6'b000000;
blue_car_bram[897] = 6'b000000;
blue_car_bram[898] = 6'b000000;
blue_car_bram[899] = 6'b000000;
blue_car_bram[900] = 6'b000000;
blue_car_bram[901] = 6'b000000;
blue_car_bram[902] = 6'b000000;
blue_car_bram[903] = 6'b000000;
blue_car_bram[904] = 6'b000000;
blue_car_bram[905] = 6'b000000;
blue_car_bram[906] = 6'b000000;
blue_car_bram[907] = 6'b000000;
blue_car_bram[908] = 6'b000000;
blue_car_bram[909] = 6'b000000;
blue_car_bram[910] = 6'b000000;
blue_car_bram[911] = 6'b000000;
blue_car_bram[912] = 6'b000000;
blue_car_bram[913] = 6'b000000;
blue_car_bram[914] = 6'b000000;
blue_car_bram[915] = 6'b000000;
blue_car_bram[916] = 6'b000000;
blue_car_bram[917] = 6'b000000;
blue_car_bram[918] = 6'b000000;
blue_car_bram[919] = 6'b000000;
blue_car_bram[920] = 6'b000000;
blue_car_bram[921] = 6'b000000;
blue_car_bram[922] = 6'b000000;
blue_car_bram[923] = 6'b000000;
blue_car_bram[924] = 6'b000000;
blue_car_bram[925] = 6'b000000;
blue_car_bram[926] = 6'b000000;
blue_car_bram[927] = 6'b000000;
blue_car_bram[928] = 6'b000000;
blue_car_bram[929] = 6'b000000;
blue_car_bram[930] = 6'b000000;
blue_car_bram[931] = 6'b000000;
blue_car_bram[932] = 6'b000000;
blue_car_bram[933] = 6'b000000;
blue_car_bram[934] = 6'b000000;
blue_car_bram[935] = 6'b000000;
blue_car_bram[936] = 6'b000000;
blue_car_bram[937] = 6'b000000;
blue_car_bram[938] = 6'b000000;
blue_car_bram[939] = 6'b000000;
blue_car_bram[940] = 6'b000000;
blue_car_bram[941] = 6'b000000;
blue_car_bram[942] = 6'b000000;
blue_car_bram[943] = 6'b000000;
blue_car_bram[944] = 6'b000000;
blue_car_bram[945] = 6'b000000;
blue_car_bram[946] = 6'b000000;
blue_car_bram[947] = 6'b000000;
blue_car_bram[948] = 6'b000000;
blue_car_bram[949] = 6'b000000;
blue_car_bram[950] = 6'b000000;
blue_car_bram[951] = 6'b000000;
blue_car_bram[952] = 6'b000000;
blue_car_bram[953] = 6'b000000;
blue_car_bram[954] = 6'b000000;
blue_car_bram[955] = 6'b000000;
blue_car_bram[956] = 6'b000000;
blue_car_bram[957] = 6'b000000;
blue_car_bram[958] = 6'b000000;
blue_car_bram[959] = 6'b000000;
blue_car_bram[960] = 6'b000000;
blue_car_bram[961] = 6'b000000;
blue_car_bram[962] = 6'b000000;
blue_car_bram[963] = 6'b000000;
blue_car_bram[964] = 6'b000000;
blue_car_bram[965] = 6'b000000;
blue_car_bram[966] = 6'b000000;
blue_car_bram[967] = 6'b000000;
blue_car_bram[968] = 6'b000000;
blue_car_bram[969] = 6'b000000;
blue_car_bram[970] = 6'b000000;
blue_car_bram[971] = 6'b000000;
blue_car_bram[972] = 6'b000000;
blue_car_bram[973] = 6'b000000;
blue_car_bram[974] = 6'b000000;
blue_car_bram[975] = 6'b000000;
blue_car_bram[976] = 6'b000000;
blue_car_bram[977] = 6'b000000;
blue_car_bram[978] = 6'b000000;
blue_car_bram[979] = 6'b000000;
blue_car_bram[980] = 6'b000000;
blue_car_bram[981] = 6'b000000;
blue_car_bram[982] = 6'b000000;
blue_car_bram[983] = 6'b000000;
blue_car_bram[984] = 6'b000000;
blue_car_bram[985] = 6'b000000;
blue_car_bram[986] = 6'b000000;
blue_car_bram[987] = 6'b000000;
blue_car_bram[988] = 6'b000000;
blue_car_bram[989] = 6'b000000;
blue_car_bram[990] = 6'b000000;
blue_car_bram[991] = 6'b000000;
blue_car_bram[992] = 6'b000000;
blue_car_bram[993] = 6'b000000;
blue_car_bram[994] = 6'b000000;
blue_car_bram[995] = 6'b000000;
blue_car_bram[996] = 6'b000000;
blue_car_bram[997] = 6'b000000;
blue_car_bram[998] = 6'b000000;
blue_car_bram[999] = 6'b000000;
blue_car_bram[1000] = 6'b000000;
blue_car_bram[1001] = 6'b000000;
blue_car_bram[1002] = 6'b000000;
blue_car_bram[1003] = 6'b000000;
blue_car_bram[1004] = 6'b000000;
blue_car_bram[1005] = 6'b000000;
blue_car_bram[1006] = 6'b000000;
blue_car_bram[1007] = 6'b000000;
blue_car_bram[1008] = 6'b000000;
blue_car_bram[1009] = 6'b000000;
blue_car_bram[1010] = 6'b000000;
blue_car_bram[1011] = 6'b000000;
blue_car_bram[1012] = 6'b000000;
blue_car_bram[1013] = 6'b000000;
blue_car_bram[1014] = 6'b000000;
blue_car_bram[1015] = 6'b000000;
blue_car_bram[1016] = 6'b000000;
blue_car_bram[1017] = 6'b000000;
blue_car_bram[1018] = 6'b000000;
blue_car_bram[1019] = 6'b000000;
blue_car_bram[1020] = 6'b000000;
blue_car_bram[1021] = 6'b000000;
blue_car_bram[1022] = 6'b000000;
blue_car_bram[1023] = 6'b000000;

    end

    // Calculate the BRAM address based on (sprite_x, sprite_y) coordinates
    wire [9:0] bram_address = (sprite_y * 32) + sprite_x;

    // Output the pixel data from the BRAM based on the address
    always @(posedge clk) begin
        pixel_data <= blue_car_bram[bram_address];
    end

endmodule