module sprite_frog (
    input [4:0] x,          // X coordinate within the sprite (0-31)
    input [4:0] y,          // Y coordinate within the sprite (0-31)
    output reg pixel        // Pixel value (1 for active, 0 for inactive)
);

    // Sprite data (32x32 binary image)
    reg [31:0] sprite_data [31:0];

    initial begin
        sprite_data[0]  = 32'b00000000000000000000000000000000;
        sprite_data[1]  = 32'b00000000000000000000000000000000;
        sprite_data[2]  = 32'b00000000000001111110000000000000;
        sprite_data[3]  = 32'b00011011000011011011000011011000;
        sprite_data[4]  = 32'b00011011000111111111100011011000;
        sprite_data[5]  = 32'b00010110001111111111110001101000;
        sprite_data[6]  = 32'b00011100011001111110011000111000;
        sprite_data[7]  = 32'b00111010010000111100001101011100;
        sprite_data[8]  = 32'b00111110110000111100001101111100;
        sprite_data[9]  = 32'b00111100111001111110011100111100;
        sprite_data[10] = 32'b00111000111111111111111100011100;
        sprite_data[11] = 32'b00111100011111111111111000111100;
        sprite_data[12] = 32'b00111111001111111111110011111100;
        sprite_data[13] = 32'b00011111101111111111110111111000;
        sprite_data[14] = 32'b00001111111110111101111111110000;
        sprite_data[15] = 32'b00000011011111111111111011000000;
        sprite_data[16] = 32'b00000001011110111101111010000000;
        sprite_data[17] = 32'b00000000111110111101111100000000;
        sprite_data[18] = 32'b00000011011110111101111011000000;
        sprite_data[19] = 32'b00000111011110111101111011100000;
        sprite_data[20] = 32'b00000111011111111111111011100000;
        sprite_data[21] = 32'b00000111011110111101111011100000;
        sprite_data[22] = 32'b00110111101110111101110111101100;
        sprite_data[23] = 32'b00110111101111111111110111101100;
        sprite_data[24] = 32'b11010111101110111101110111101011;
        sprite_data[25] = 32'b11111011110111111111101111011111;
        sprite_data[26] = 32'b01111101110111111111101110111110;
        sprite_data[27] = 32'b11111111110001111110001111111111;
        sprite_data[28] = 32'b11111111100000011000000111111111;
        sprite_data[29] = 32'b00111111100000000000000111111100;
        sprite_data[30] = 32'b00000110000000000000000001100000;
        sprite_data[31] = 32'b00000000000000000000000000000000;
    end

    // Output the pixel value based on the (x, y) coordinates
    always @(*) begin
        pixel = sprite_data[y][x];
    end

endmodule
